{
"##0_entertainment_access##":"Denna boning har inte tillgång till underhållning överhuvudtaget"
"##1_entertainment_access##":"Denna boning har knappt tillgång till underhållning"
"##2_entertainment_access##":"Denna boning har viss tillgång till underhållning"
"##3_entertainment_access##":"Denna boning har mycket begränsad tillgång till underhållning"
"##4_entertainment_access##":"Denna boning har rimlig tillgång till underhållning"
"##5_entertainment_access##":"Denna boning har begränsad tillgång till underhållning"
"##6_entertainment_access##":"Denna boning har god tillgång till underhållning"
"##7_entertainment_access##":"Denna boning har mycket god tillgång till underhållning"
"##8_entertainment_access##":"Denna boning har utmärkt tillgång till underhållning"
"##9_entertainment_access##":"Denna boning har tillgång till all underhållning som kan önskas"
"##academies##":"Högskolor"
"##academy_full_work##":"Denna högskola används, och ungdomarna i stadsdelen lär sig sociala färdigheter."
"##academy_info##":"En del ungdomar som går ut skolorna går vidare och studerar avancerad retorik och historia vid högskolan. Alla kulturella medborgare har en akademisk bakgrund."
"##academy_no_workers##":"Denna högskola används inte, och är därför värdelös för lokalsamhället."
"##academy_trained##":"Utbildad på högskola"
"##academy##":"Högskola"
"##accept_deity_status##":"Acceptera ställningen som kejsare!"
"##accept_goods##":"Acceptera varor"
"##accept_promotion##":"Acceptera befordran"
"##accept##":"Acceptera"
"##accepting##":"Accepterar"
"##access_ramp##":"Åtkomstramp"
"##actor_average_life##":"Livet här är helt enkelt ljuvligt."
"##actor_gods_angry##":"Aaagh!! Gudarna är vreda. Vi går under!"
"##actor_good_life##":"Den här staden är inte så illa."
"##actor_high_workless##":"Det är så stor arbetslöshet att jag inte förmår lära mig mina repliker."
"##actor_low_entertainment##":"Jag arbetar så hårt jag förmår, men underhållningen i staden räcker inte till på långa vägar."
"##actor_need_workers##":"Det finns helt enkelt inte tillräckligt med arbetare i staden."
"##actor_so_hungry##":"Jag kan inte uppträda utan mer mat."
"##actor##":"Skådespelare"
"##actorColony_bad_work##":"Jag har ingen personal utöver mig själv. Jag kan inte arbeta under dessa förhållanden! Som bäst kan jag utbilda en skådespelare på tre månader."
"##actorColony_full_work##":"Det är med nöje vi tillkännager att vi, med full sysselsättning, kan hjälpa upp till fyra nya skådespelare varje månad."
"##actorColony_need_some_workers##":"Vi är något underbemannade, och kan därför endast utbilda två nya skådespelare per månad."
"##actorColony_no_workers##":"Denna koloni är övergiven. Utan tillgång till mentorer kan inga nya skådespelare utbildas."
"##actorColony_patrly_workers##":"Vi har bara halva personalstyrkan, och kan därför endast utbilda en skådespelare under nästa månad."
"##actorColony_slow_work##":"Vi lider av svår personalbrist, och kommer att få kämpa för att utbilda en ny skådespelare under de kommande två månaderna."
"##actorColony##":"Skådespelarkoloni"
"##ad##":"eKr"
"##adjust_exact##":"Ställ in den exakta summa du vill donera"
"##adjust_tax_rate##":"Justera skattenivån i staden"
"##administration_building##":"Administrativa- och regeringsbyggnader"
"##advanced_houseinfo##":"Avancerad information om detta hus"
"##advchief_crime##":"Brott"
"##advchief_education##":"Utbildning"
"##advchief_employers_ok##":"Staden har inga sysselsättningsproblem"
"##advchief_employment##":"Arbete"
"##advchief_finance##":"Finanser"
"##advchief_food_consumption##":"Matförbrukning"
"##advchief_food_stocks##":"Matförråd"
"##advchief_havedeficit##":"Tillgångarna har i år minskat med"
"##advchief_haveprofit## ":"Tillgångarna har i år stigit med"
"##advchief_health_awesome_clinic##":"Stadens hälsosituation är utmärkt, inga väntetider alls för besök till lokala läkare."
"##advchief_health_awesome##":"Stadens hälsosituation är utmärkt"
"##advchief_health_bad_clinic##":"Stadens hälsosituation är dålig, dina överansträngda läkare fruktar en dödlig epidemi."
"##advchief_health_bad##":"Stadens hälsosituation är dålig"
"##advchief_health_good_clinic##":"Stadens hälsosituation är nästan perfekt, läkarnas kliniker är nästan tomma."
"##advchief_health_good##":"Stadens hälsosituation är nästan perfekt"
"##advchief_health_high_clinic##":"Stadens hälsosituation är bra, dina medborgare lider bara av enklare sjukdomar."
"##advchief_health_high##":"Stadens hälsosituation är bra"
"##advchief_health_less_clinic##":"Stadens hälsosituation är dålig, mat och kliniker skulle förbättra hälsan."
"##advchief_health_less##":"Stadens hälsosituation är ganska dålig"
"##advchief_health_low##":"Stadens hälsosituation är förfärande"
"##advchief_health_lower##":"Stadens hälsosituation är förfärande, pest kommer med all säkerhet bryta ut."
"##advchief_health_middle_clinic##":"Stadens hälsosituation är tillfredsställande, klinikerna håller farliga epidemier borta."
"##advchief_health_middle##":"Stadens hälsosituation är tillfredsställande"
"##advchief_health_perfect_clinic##":"Stadens hälsosituation är perfekt, dina tomma kliniker utgör ett exempel genom hela imperiet."
"##advchief_health_perfect##":"Stadens hälsosituation är perfekt"
"##advchief_health_simple_clinic##":"Stadens hälsosituation är mindre bra"
"##advchief_health_simple##":"Stadens hälsosituation är inte bra, se till att dina medborgare har mat och kliniker."
"##advchief_health_terrible_clinic##":"Stadens hälsosituation är fruktansvärd, klinikerna hinner inte med, sjukdomar är nästan oundvikliga."
"##advchief_health_terrible##":"Stadens hälsosituation är fruktansvärd"
"##advchief_health_verygood_clinic##":"Stadens hälsosituation är mycket bra, medborgarnas småkrämpor hanteras snabbt av lokala läkare."
"##advchief_health_verygood##":"Stadens hälsosituation är mycket bra"
"##advchief_health##":"Hälsa"
"##advchief_high_crime_in_district##":"Vissa områden har hög kriminalitet"
"##advchief_high_crime##":"Stor kriminalitet råder i staden"
"##advchief_low_crime##":"Det finns lite brottslighet här, ingenting allvarligt."
"##advchief_military##":"Militär"
"##advchief_needworkers##":"Staden saknar"
"##advchief_sentiment##":"Stämning"
"##advchief_some_need_academy##":"Vissa medborgare vill ha fler skolor"
"##advchief_some_need_barber##":"Vissa medborgare behöver barberare"
"##advchief_some_need_baths##":"Vissa medborgare behöver badhus"
"##advchief_some_need_doctors##":"Vissa medborgare behöver läkarkliniker"
"##advchief_some_need_education##":"Medborgarna kräver mer utbildning"
"##advchief_some_need_hospital##":"Vissa medborgare behöver sjukhus"
"##advchief_some_need_library##":"Vissa medborgare vill ha fler bibliotek"
"##advchief_which_crime_in_district##":"Vissa områden har mindre problem"
"##advchief_which_crime##":"Brottsligheten håller på att bli ett problem."
"##advchief_workless##":"Staden har en arbetslöshet på"
"##adve_administration_religion##":"Styrelse/Religion"
"##adve_engineers##":"Konstruktion"
"##adve_entertainment##":"Underhållning"
"##adve_food##":"Livsmedelsproduktion"
"##adve_health_education##":"Hälsa och utbildning"
"##adve_industry_and_trade##":"Industri och handel"
"##adve_military##":"Militär"
"##adve_prefectures##":"Prefekturer"
"##adve_water##":"Vattenförsörjning"
"##advemp_emperor_favour##":"Popularitet"
"##advemployer_panel_denaries##":""
"##advemployer_panel_haveworkers##":""
"##advemployer_panel_needworkers##":""
"##advemployer_panel_priority##":""
"##advemployer_panel_romepay##":"Rom betalar"
"##advemployer_panel_salary##":"Löner"
"##advemployer_panel_sector##":""
"##advemployer_panel_title##":"Arbetstilldelning"
"##advemployer_panel_workers##":""
"##advemployer_panel_workless##":"Arbetslös arbetsstyrka "
"##advice_at_culture##":"Klicka här för information om din kulturställning"
"##advisors##":"Senat"
"##advlegion_noalarm##":"Vi har inga rapporter om hot mot staden"
"##advlegion_norequest##":"Vi har inte fått någon begäran om hjälp från imperiet"
"##advlegion_window_title##":"Legionstatus"
"##advpopulation_text_census##":"Befolkningssammansättning efter ålder (år)"
"##advpopulation_text_society##":"Befolkningssammansättning efter inkomst"
"##advpopulation_title_census##":"Befolkning - Folkräkning"
"##advpopulation_title_population##":"Befolkning - Historia"
"##advpopulation_title_society##":"Befolkning - Samhälle"
"##aedile##":"Edil"
"##age_ad##":"eKr"
"##age_bc##":""
"##also_fountain_in_well_area##":"Denna brunn är överflödig för tillfället, eftersom alla hus som den betjänar tar sitt vatten från en fontän."
"##amazing_prosperity_this_city##":"Det fantastiska välståndet i den här staden är det stora samtalsämnet i Rom!"
"##amphitheater_full_work##":"Denna amfiteater erbjuder sitt samhälle både intressant gladiatorkamp och pjäser med lokala skådespelare."
"##amphitheater_have_never_show##":"Denna amfiteater har sällan några föreställningar. Den behöver skådespelare och gladiatorer."
"##amphitheater_have_only_battles##":"Denna amfiteater erbjuder gladiatorkamp som förströelse. Den söker skådespelare för att sätta upp några pjäser."
"##amphitheater_have_only_shows##":"Denna amfiteater sätter upp pjäser med lokala aktörer. Den kan attrahera större publik om den även har gladiatorer."
"##amphitheater_haveno_gladiator_bouts##":"Ingen gladiatorkamp för närvarande"
"##amphitheater_haveno_shows##":"Inga pjäser för närvarande"
"##amphitheater_no_access##":"Detta hus har inte tillgång till en amfiteater"
"##amphitheater_no_workers##":"Denna amfiteater är stängd. Den har inga anställda, och erbjuder ingen förströelse åt det lokala samhället."
"##amphitheater##":"Amfiteater"
"##amphitheatres##":"Amfiteatrar"
"##angry##":"Arga"
"##animal_contests_run##":"Djurtävlingarna pågår ytterligare"
"##aqueduct_info##":"Akvedukter gör det möjligt att konstruera reservoarer långt från vatten, vilket gör det möjligt för fontäner att förse staden med vatten."
"##aqueduct_no_water##":"Denna akvedukt transporterar inte vatten mellan reservoarer eftersom den saknar vattenkälla."
"##aqueduct_work##":"Denna akvedukt transporterar vatten mellan reservoarer."
"##aqueduct##":"Akvedukt"
"##arabian_stallions##":"Arabiska hingstar"
"##architect_salary##":"Arkitektlön på"
"##architect##":"Arkitekt"
"##army_marker##":"Armémarkör"
"##arrange_festiable_for_this_god##":"Arrangera en festival till denna guds ära"
"##arrow##":"Pil"
"##averange_crime_risk##":"Detta är ett område med hög brottslighet. De boende är missnöjda, och gatorna är farliga"
"##avesome_amphitheater_access##":"Detta hus passerades nyligen av en gladiator. Det kommer att ha tillgång till amfiteater under lång tid framåt"
"##avesome_clinic_access##":"Detta hus passerades nyligen av en läkare. Det kommer att ha tillgång till en klinik under lång tid framåt"
"##avesome_college_access##":"Detta hus passerades nyligen av en lärare. Det kommer att ha tillgång till högskola under lång tid framåt"
"##avesome_colloseum_access##":"Detta hus passerades nyligen av en lejontämjare. Det kommer att ha tillgång till ett colosseum under lång tid framåt"
"##avesome_hippodrome_access##":"Detta hus har nyligen passerats av en körsven. Det kommer att ha tillgång till hippodrom under lång tid framåt"
"##avesome_hospital_access##":"Detta hus passerades nyligen av en kirurg. Det kommer att ha tillgång till sjukhus under lång tid framåt"
"##avesome_library_access##":"Detta hus har nyligen passerats av en bibliotekarie. Det kommer att ha tillgång till bibliotek under lång tid framåt"
"##avesome_school_access##":"Detta hus passerades nyligen av ett skolbarn. Det kommer att ha tillgång till skola under lång tid framåt"
"##avesome_theater_access##":"Detta hus passerades nyligen av en skådespelare. Det kommer att ha tillgång till teater under lång tid framåt"
"##awesome_amphitheater_access##":"Detta hus har tillgång till amfiteater"
"##awesome_barber_access##":"Detta hus har tillgång till barberare"
"##awesome_barber_access##":"Detta hus passerades nyligen av en barberare. Det kommer att ha tillgång till en barberare under lång tid framåt"
"##awesome_baths_access##":"Detta hus har tillgång till badhus"
"##awesome_baths_access##":"Detta hus passerades nyligen av en badhusarbetare. Det kommer att ha tillgång till badhus under lång tid framöver"
"##awesome_colloseum_access##":"Detta hus har tillgång till colosseum"
"##awesome_doctor_access##":"Detta hus har tillgång till en klinik"
"##awesome_entertainment_access##":"Denna boning har tillgång till flera platser för underhållning"
"##bad_house_quality##":"Den totala kvaliteten på byggnaderna i din stad inverkar negativt på denna ställning."
"##balance##":"Balans"
"##ballista##":"Kastmaskin"
"##barbarian_attack_text##":""
"##barbarian_attack_title##":"Fiender attackerar staden"
"##barbarian_warrior##":"En barbarisk soldat"
"##barber_access##":"Barberartillgång"
"##barber_average_life##":"Är inte den här staden ett riktigt klipp?"
"##barber_full_work##":"Denna barberarlokal används, och ortsbefolkningen är vältrimmad."
"##barber_gods_angry##":"Gudarna är vreda. Jag önskar att ståthållaren skulle bygga fler tempel."
"##barber_good_life##":"Rakning eller klippning, medborgare? Livet här är lätt att leva, inte sant?"
"##barber_high_workless##":"Arbetslösheten är så hög att den får håret att stå på ända!"
"##barber_info##":"Ingen civiliserad man visar sig orakad offentligt! Alla medborgare behöver regelbundet besöka en barberare för att kunna avancera i samhället."
"##barber_need_colloseum##":"Efter en dag med rakning och klippning vill jag se en trevlig lejonstrid. Men det går inte att uppbringa här."
"##barber_need_workers##":"Det saknas många arbetare här."
"##barber_no_access##":"Detta hus har inte tillgång till en barberare"
"##barber_no_workers##":"Denna barberarlokal används inte, och är därför värdelös för lokalsamhället."
"##barber_shop##":"Barberare"
"##barber_so_hungry##":"En hårklippning får dig att glömma hungern. Och det är många hungriga i den här staden."
"##barber##":"Barberare"
"##barbers##":"Barberare"
"##barracks_bad_weapons_bad_workers##":"Med minimipersonal och inga vapenupplag får vi kämpa för att utbilda till och med de mest enkla trupper."
"##barracks_bad_weapons_need_some_workers##":"Vi saknar några anställda och utbildar soldater långsammare än vanligt. Utan vapenupplag kan vi inte utbilda några nya legionärer."
"##barracks_bad_weapons_slow_workers##":"Vi är underbemannade och saknar vapen, vi kan bara långsamt utbilda stödtrupper."
"##barracks_city_not_need_soldiers##":"Vi utbildar för närvarande inga rekryter eftersom vi inte har fått någon begäran från stadens fort eller torn om nya styrkor."
"##barracks_full_work##":"Vi utbildar nya soldater med maximal effektivitet och vi har vapen för att utbilda alla typer av soldater."
"##barracks_have_weapons_bad_workers##":"Med minimipersonal utbildar vi nya soldater mycket långsamt trots att vi har de vapen som krävs för att utbilda alla typer av soldater."
"##barracks_have_weapons_slow_workers##":"Vi är underbemannade och utbildar nya soldater långsamt, men vi har de vapen som krävs för att utbilda alla typer av soldater."
"##barracks_info##":"Ingen kan gå med i en romersk legion utan att först komma hit. Alla nya rekryter kommer hit."
"##barracks_need_some_workers##":"Pga. personalbrist utbildar vi nya soldater långsammare än vanligt men vi har de vapen som krävs för att utbilda alla typer av soldater."
"##barracks_no_weapons##":"Vi kan utbilda stödtrupper mycket snabbt, men utan vapenupplag kan vi inte utbilda några nya legionärer."
"##barracks##":"Förläggningar"
"##bath_1##":"Badhus"
"##bath_access##":"Badtillgång"
"##bath_no_access##":"Detta hus har inte tillgång till ett fungerande badhus"
"##bath##":"Badhus"
"##bathlady_so_hungry##":"Folk har inte ätit på så länge att deras revben börjar sticka ut, vilket syns på badhuset."
"##bathlady##":"Badarbetare"
"##baths_full_work##":"Detta badhus används, besökarna blir rena och avslappnade."
"##baths_info##":"Civiliserade människor badar minst en gång om dagen. Utöver bättre hälsa utgör baden även en önskvärd träffpunkt med olika rekreativa aktiviteter."
"##baths_need_reservoir##":"Detta badhus behöver en rörledning till en reservoar."
"##baths_no_workers##":"Detta badhus används inte, och är därför värdelöst för lokalsamhället."
"##baths##":"Badhus"
"##bc##":"fKr"
"##beatifull_villa##":"Stor villa"
"##beatyfull_insula##":"Storslagen Insulae"
"##become_trade_center##":"Utse till handelscentral"
"##below_average##":"Under medel"
"##better_class_road##":"En finare typ av väg"
"##big_domus##":"Stor Insula"
"##big_hovel##":"Stort skjul"
"##big_hut##":"Stort hus"
"##big_palace##":"Stort palats"
"##big_shack##":"Stor koja"
"##big_tent##":"Stor tält"
"##big_villa##":"Stor villa"
"##bldm_factory##":"Verkstäder"
"##bldm_farm##":"Jordbruk"
"##bldm_raw_materials##":"Råmaterial"
"##bldm_raw##":"Råmaterial"
"##bolt##":"Armborst"
"##bridge_extends_city_area##":"Denna bro ger oss mer mark, men ger fri passage både för medborgare och fiender!"
"##bridge##":"Bro"
"##bridges##":"Broar"
"##briton##":"En britt"
"##britons##":"Britter"
"##broke_empiretax_warning##":"Din oförmåga att betala tribut till Rom utmålar din stad som misslyckad."
"##broke_empiretax_with2years_warning##":"Din fortsatta oförmåga att lämna tribut till Rom skadar ditt rykte."
"##btn_showprice_tooltip##":"Visar import-/exportpriser för alla varor, som anbefallt av Rom"
"##build_fishing_boat##":"Vi bygger båtar på beställning från en fiskehamn i staden."
"##build_housing##":"Bygg bostäder"
"##build_markets_to_distribute_food##":"Bygg marknader för att distribuera maten som lagrats här"
"##build_road_tlp##":"Bygg vägar"
"##building_need_road_access##":""
"##buildings##":"Byggnation"
"##burning_ruins##":"Brinnande ruin"
"##buy_price##":"Köparna betalar"
"##caesar_assign_new_title##":"Caesar har befordrat dig till graden"
"##caesar_salary##":"Caesars lön på"
"##caesarea_win_text##":"Så Caesareas förre ståthållare ska alltså få behålla livet? Att rädda staden ur krisen är verkligen en bedrift. Jag kanske ska låta dig välja vilket land vi ska utvisa honom till."
"##can_build_only_one_of_building##":"Du kan endast ha en byggnad av denna typ"
"##cancel##":"Avbryt"
"##cancelBtnTooltip##":"Avbryt denna operation"
"##cant_calc_prosperity##":"Din stad är ny. Vi har inte haft möjlighet att bedöma ditt välstånd än!"
"##cant_demolish_bridge_with_people##":"Kan inte förstöra bro med människor på"
"##captured_city##":"En erövrad stad"
"##carthaginian_soldier##":"En karthagisk soldat"
"##carthago_win_text##":"Tack vare din briljanta insats ligger det karthagiska hotet äntligen bakom oss. Våra forna fiender är nu laglydiga romerska medborgare. I alla fall de som ännu är i livet!"
"##cartPusher_average_life##":"...knappast roligt, men att få bo i denna fina stad gör det mödan värt."
"##cartPusher_cantfind_destination##":"Det skulle gå snabbare att dra varorna till Rom än dit jag ska."
"##cartPusher_gods_angry##":"...religiös, men inte ens jag skulle behandla gudarna på det här sättet."
"##cartPusher_good_life##":"Stad som stad... Den här verkar rätt bra."
"##cartPusher_high_workless##":"...min fru har slutat tjata om att jag ska skaffa mig ett nytt arbete."
"##cartPusher_low_entertainment##":"...vagnar. Det är mer underhållande än resten av den här staden."
"##cartPusher_need_workers##":"Vart man än kommer i staden finns det lediga arbeten."
"##cartPusher_so_hungry##":"...dagen kräver styrka. Hur ska en vagndragare kunna arbeta utan mat?"
"##ceres_badmood_info##":"Ceres missnöje är farligt, eftersom hon skyddar folket från dåliga skördar och hungersnöd."
"##ceres_desc##":"Jordbruk"
"##ceres_goodmood_info##":"Ceres skänker fruktsamhet åt jorden, och får plantorna att växa. Blidka henne, eller bered dig på hungersnöd."
"##changesalary_greater_salary##":"Varning: Betala dig själv en lön som överstiger din grad imponerar inte på kejsaren."
"##charioteer_school_full_work##":"Det är med nöje vi tillkännager att vi, med full sysselsättning, kan slutföra upp till fyra nya vagnar varje månad."
"##charioteer_school_need_some_workers##":"Vi är något underbemannade, och kan därför endast tillverka två nya vagnar per månad."
"##charioteer_school_patrly_workers##":"Vi har bara halva personalstyrkan, och kan därför endast tillverka en vagn under nästa månad."
"##charioteer##":"Körsven"
"##charioter_so_hungry##":"Hungrig? Jag kan äta en häst, så lite mat finns det."
"##chatioteer_school_bad_work##":"Jag har ingen personal utöver mig själv. Jag kan inte arbeta under dessa förhållanden! Jag kan bara bygga en vagn på tre månader."
"##chatioteer_school_info##":"De hantverkare som arbetar här bygger snabba, kraftiga vagnar och utbildar förarna. Kapplöpningarna i hippodromen är mycket populära."
"##chatioteer_school_no_workers##":"Utan hantverkare kan inga nya vagnar produceras. Som resultat kan hippodromen, om den är i drift, bli lidande."
"##chatioteer_school_slow_work##":"Vi lider av svår personalbrist, och kommer att få kämpa för att bygga en enda ny vagn under de kommande två månaderna."
"##chatioteer_school##":"Skola för körsvenner"
"##chief_advisor##":"Huvudrådgivare"
"##children##":"Barn"
"##citizen_are_rioting##":"Medborgarna gör uppror!"
"##citizen_gods_angry##":"Detta är en hednisk stad. Den behöver fler tempel."
"##citizen_gods_angry3##":"Den här ståthållaren har ingen respekt för gudarna."
"##citizen_good_education##":"Den här staden är mer kultiverad än någon annan i riket!"
"##citizen_high_workless10##":"Arbetslösheten är så hög att hela staden mår dåligt."
"##citizen_high_workless2##":"Om jag inte får arbete snart, måste jag flytta till en annan stad."
"##citizen_high_workless4##":"Jag har aldrig sett så många arbetslösa medborgare förut."
"##citizen_low_entertainment4##":"Man kan inte roa sig alls på det här stället."
"##citizen_low_salary##":"Min hund skulle inte arbeta för de löner de betalar här. Jag ger mig av."
"##citizen_need_workers3##":"Staden lider stor brist på arbetare."
"##citizen_need_workers5##":"Staden behöver fler arbetare!"
"##citizen_salary##":"Medborgarlön på"
"##citizen##":"Medborgare"
"##citizens_additional_rooms_for##":"Extra utrymme för"
"##city_cyrene##":"Cyrene"
"##city_damascus##":"Damascus"
"##city_fire_text##":"Prefekterna kunde inte nå hit i tid för att rädda byggnaden. När elden har brunnit ut kommer endast spillror att finnas kvar på denna plats."
"##city_fire_title##":""
"##city_has_debt##":"Staden har en skuld till Rom på"
"##city_has_runout_debt##":""
"##city_have_goods_for_request##":""
"##city_have##":"Stadens skattkammare har tillgångar på"
"##city_health##":"Hälsosituation"
"##city_loathed_you##":"Du föraktas i hela staden"
"##city_need_more_workers##":"Din stad kräver fler arbetare"
"##city_sounds_off##":"Stadsljud är AV"
"##city_sounds_on##":"Stadsljud är PÅ"
"##city##":"Stad"
"##citychart_census##":"Folkräkning"
"##citychart_population##":"Historia"
"##citychart_society##":"Samhälle"
"##clay_factory_stock##":"Lagrad lera,"
"##clay_pit_bad_work##":"Det finns nästan inga som gräver vid detta lertag, och produktionen står nästan still. Mycket lite lera produceras under det kommande året."
"##clay_pit_full_work##":"Detta lertag har alla anställda det behöver, och arbetar fullt ut med att producera lera."
"##clay_pit_info##":"Tag lera och handla med, eller leverera den till krukmakerier. Folket behöver krukor för att bebo Insulaen."
"##clay_pit_need_close_to_water##":"Bygg lertag nära vattnet"
"##clay_pit_need_some_workers##":"Detta lertag utnyttjar inte full kapacitet. Som resultat kommer lerproduktionen att gå något långsammare."
"##clay_pit_no_workers##":"Detta lertag har inga anställda. Produktionen har upphört."
"##clay_pit_patrly_workers##":"Detta lertag är underbemannat, och det tar längre tid att producera leran än vad det borde."
"##clay_pit_patrly_workers##":"Detta brott är underbemannat, och det tar längre tid än det borde att producera marmorn."
"##clay_pit##":"Lertag"
"##clay##":"Lera"
"##clear_land_caption##":"Tomt land"
"##clear_land_text##":"Detta landområde kan byggas på efter behov. Det ger fri passage både åt egna soldater och åt fiendesoldater."
"##clear_land##":"Röj marken"
"##clerk_salary##":"Bokhållarlön på"
"##clerk##":"Bokhållare"
"##click_here_that_stacking##":"Klicka här för att hamstra"
"##click_here_that_use_it##":"Klicka här för att stänga av hamstring"
"##click_item_for_start_trade##":"Klicka på en vara"
"##click_on_city_for_info##":"Klicka på en stad för att få information"
"##clinic_full_work##":"Denna klinik används, och betjänar lokalsamhället."
"##clinic_info##":"Läkares förbättrar medborgarnas hälsa genom sina hembesök i de stadsdelar som ingår i deras runda. Blomstrande områden vill ha en klinik."
"##clinic_no_workers##":"Denna klinik används inte, och är därför värdelös för lokalsamhället."
"##clinic##":"Klinik"
"##clinics##":"Kliniker"
"##colege_access_perfectly##":"Områden som kräver utbildningsmöjligheter har tillgång till dem, men fler högskolor skulle minska storleken på klasserna."
"##collapse_available_damage_risk##":"Mycket stor risk för kollaps"
"##collapse_immitent##":"Överhängande risk för kollaps"
"##collapsed_ruins_info##":"Dessa spillror av gamla byggnader gör marken mindre åtråvärd."
"##colloseum_haveno_animal_bouts##":"Inga djurkamper för närvarande"
"##colloseum_haveno_gladiator_bouts##":"Ingen aktuell gladiatorkamp"
"##colloseum_haveno_gladiatorpit##":"Bygg en gladiatorskola för att arrangera matcher här"
"##colloseum_info##":"Colosseum och amfiteatrar behöver alltid nya gladiatorer för att ersätta förlorarna."
"##colloseum_no_workers##":"Detta colosseum är stängt. Utan anställda är det värdelöst som rekreationsanläggning."
"##colloseum##":"Colosseum"
"##colloseums##":"Colosseum"
"##colosseum_no_access##":"Detta hus har ingen tillgång till ett colosseum"
"##column_info##":"Kolonnformation"
"##comerceBtnTooltip##":""
"##commerce##":"Handel"
"##congratulations##":"Gratulerar"
"##consul_salary##":"Konsulslön på"
"##consul##":"Konsul"
"##contaminted_water##":"Förorenat vatten"
"##continue##":""
"##corinthus##":"Corinthus"
"##cost_2_open##":"Kostnad att öppna"
"##cost##":"Kostnad"
"##costs##":"kostnader"
"##coverage##":"Täckning i staden"
"##crack##":"Spricka"
"##credit##":"Utgifter"
"##current_game_speed_is##":""
"##current_year_notpay_tribute_warning##":"Du har inte betalat tribut detta året. Spara lite pengar i din skattkammare så att du kan göra din årliga betalning."
"##cursed_by_mars##":"Förbannad av Mars!"
"##damage##":"Skador"
"##damascus_somewhat_dangerous_province##":"Damaskus: en relativt farlig provins"
"##damascus_win_text##":"Ännu en gång har du uppnått vad svagare män kallar omöjligt. Hela östern åsåg din balansgång i Damaskus. Nu kan jag tryggt hämta hem några av mina syriska legioner."
"##dangerous_crime_risk##":"Detta område är farligt."
"##date_tooltip##":""
"##date##":"Datum"
"##day_longer_in_that_tent##":"En dag till i det tältet och jag hade exploderat"
"##day##":"Dag"
"##days##":"Dagar"
"##debet##":"Inkomst"
"##dedicate_fectival_ceres##":"Tillägna Ceres en festival"
"##dedicate_fectival_mars##":"Tillägna Mars en festival"
"##dedicate_fectival_mercury##":"Tillägna Merkurius en festival"
"##dedicate_fectival_neptune##":"Tillägna Neptunus en festival"
"##dedicate_fectival_venus##":"Tillägna Venus en festival"
"##defensive_formation_text##":"En mycket defensiv formation. Nästan omöjlig att penetreras av missiler."
"##delete_game##":""
"##delete_object##":"Radera objekt"
"##delete_this_message##":"Radera detta meddelande"
"##delighted##":"Förtjusta"
"##deliver##":"Hämta varor"
"##delivery_boy##":"Springpojke"
"##demand##":"Krav"
"##demands_3_religion##":"Krav på tillgång till en tredje religion"
"##denarii_short##":""
"##desirability_indiffirent_area##":"Dina medborgare ser varken positivt eller negativt på detta område"
"##desirability_pretty_area##":"Detta land är ett eftertraktat område, vad gäller dina medborgare"
"##desirability##":"Önskvärdhet"
"##destroy_bridge_warning##":"Sätt tillbaka Caesar III CD'n i CD-ROM enheten"
"##destroy_bridge##":"CD saknas"
"##destroy_fort##":"Förstör ett fort"
"##devastate_granary##":"Töm sädesmagasin"
"##devastate_warehouse##":"BÖRJA tömma magasin"
"##developers##":""
"##difficulty##":""
"##disasterBtnTooltip##":""
"##dispatch_force##":"Sänd iväg undsättningsstyrka?"
"##dispatch_gift##":"Sänd en gåva"
"##dispatch_git_title##":"Sänd gåva till kejsaren"
"##dispatch_goods?##":"Sända iväg varor?"
"##distant_city##":"En avlägsen stad"
"##distribution_center##":"Distributionscentral"
"##dn_collected_this_year##":"denarer har betalats hittills i år"
"##dn_for_open_trade##":"för att öppna handelsväg"
"##dn_per_month##":"denarer per månad"
"##dn's##":"Avsluta byggare"
"##dn##":"Spara karta"
"##dock_bad_work##":"Vi har mycket få hamnarbetare så det kommer att ta lång tid att lasta och lossa de fartyg som anlöper hamnen."
"##dock_bad_work##":"Vi kan inte betjäna det förtöjda fartyget utan hamnarbetare!"
"##dock_busy_bad_work##":"Vi betjänar det förtöjda fartyget, men har för få hamnarbetare, detta kommer att ta tid."
"##dock_busy_patrly_workers##":"Vi betjänar det förtöjda fartyget, trots att vi inte har tillräckligt med anställda, så det kommer att ta längre tid än det borde."
"##dock_cart_returning_from":"Vår vagn återvänder från en leverans."
"##dock_cart_taking_goods##":"Vår vagn för varorna till annan plats."
"##dock_cart_wait##":"Vår vagn är här och väntar på nya order."
"##dock_full_work##":"Vi har full arbetsstyrka och kommer att kunna lasta och lossa inkommande fartyg."
"##dock_info##":"Hamnarbetarna hämtar varor som vi köper från lagerlokalen."
"##dock_info##":"Handelsskepp från hela riket lägger till här för att leverera importvaror och hämta exportvaror. Du kan inte bedriva sjöhandel utan en handelshamn."
"##dock_need_some_workers##":"Vi är underbemannade och därför kommer det att ta lite längre tid än vanligt att lasta och lossa de fartyg som anlöper hamnen."
"##dock_no_workers##":"Vi har inga hamnarbetare och kan därför inte lasta eller lossa några fartyg som kommer till hamnen."
"##dock##":"Handelshamn"
"##docked_buying_selling_goods##":"Ligger vid kaj, köper och säljer varor"
"##doctor_average_life##":"Detta är en fantastisk stad."
"##doctor_gods_angry##":"Gudarna är upprörda. Om vi inte respekterar dem, kommer vi att få känna på deras vrede."
"##doctor_good_life##":"Stadens invånare tycks vara vid god hälsa."
"##doctor_high_workless##":"Arbetslösheten är mycket hög. Jag funderar på att ge mig av."
"##doctor_low_entertainment##":"Staden är så trist att mina patienter frågar om jag kan bota kronisk uttråkning!"
"##doctor_need_workers##":"Var hälsad! Det saknas många arbetare här."
"##doctor_no_access##":"Detta hus har inte tillgång till en klinik"
"##doctor_so_hungry##":"Folk är undernärda, men det saknas mat att bota det med."
"##donation_is##":"Donationen är"
"##donations##":"Donerat"
"##donationwnd_exit_tip##":"Lämna donationsskärmen"
"##donot_organize_festival##":"Organisera ingen festival"
"##east##":"Öst"
"##edadv_need_better_access_school_or_colege##":"Bättre skola eller högskola och tillgång till bibliotek skulle förbättra vissa områden i staden. Man skall inte behöva gå långt för att lära sig något!"
"##edil_salary##":"Edillön på"
"##education_advisor_title##":"Utbildning"
"##education_awesome##":"Alla som kräver utbildningsmöjligheter i staden har dem, och dessa är perfekta i hela staden."
"##education_full_access##":"Detta hus har tillgång till skola, bibliotek och högskola"
"##education_have_academy_access##":"Detta hus har tillgång till högskola"
"##education_have_no_access##":"Detta hus har ingen grundläggande tillgång till skolor eller bibliotek"
"##education_have_school_library_access##":"Detta hus har tillgång till skola och bibliotek"
"##education_have_school_or_library_access##":"Detta hus har tillgång till skola eller bibliotek"
"##education_objects##":"Utbildningsbyggnader"
"##education##":"Utbildning"
"##educationBtnTooltip##":""
"##egift_chest_of_sapphire##":"En kista med safirer"
"##egift_educated_slave##":"En utbildad slav"
"##egift_egyptian_glassware##":"Egyptiska glasvaror"
"##egift_gaulish_bodyguards##":"Galliska livvakter"
"##egift_generous##":"Generös:"
"##egift_gepards_and_giraffes##":"Geparder och giraffer"
"##egift_golden_chariot##":"En gyllene vagn"
"##egift_gree_manuscript##":"Ett grekiskt manuskript"
"##egift_lavish##":"Frikostig:"
"##egift_modest##":"Blygsam:"
"##egift_persian_carpets##":"Persiska mattor"
"##egift_soldier_from_pergamaum##":"En soldat från Pergamon"
"##egift_troupe_preforming_slaves##":"En grupp uppträdande slavar"
"##emigrant_high_workless##":"Vet ni var det kan finnas arbete? Jag måste få ett arbete."
"##emigrant_no_home##":"Jag har ingenstans att bo."
"##emigrant_no_work_for_me##":"Jag har fått nog av detta ställe. Det finns inget arbete här."
"##emigrant_thrown_from_house##":"Jag har blivit utkastad från mitt hem!"
"##emigrant##":"Emigrant"
"##empbutton_low_work##":"Fungerar dåligt. Tilldela fler människor till vår sektor"
"##empbutton_simple_work##":"Fungerar, men fler arbetare skulle kunna tilldelas oss"
"##empbutton_tooltip##":"Klicka här för att fastställa en prioritet för denna arbetskraftskategori"
"##emperor_favour_00##":"Kejsaren är rasande på dig."
"##emperor_favour_01##":"Kejsaren är så otroligt arg att han talar om att landsförvisa dig."
"##emperor_favour_02##":"Kejsaren är vansinnigt arg på dig."
"##emperor_favour_03##":"Kejsaren är mycket arg på dig."
"##emperor_favour_04##":"Kejsaren är arg på dig."
"##emperor_favour_05##":"Kejsaren är extremt missnöjd med dig."
"##emperor_favour_06##":"Kejsaren är mycket missnöjd med dig."
"##emperor_favour_07##":"Kejsaren är missnöjd med dig."
"##emperor_favour_08##":"Kejsaren är något missnöjd med dig."
"##emperor_favour_09##":"Kejsaren är tveksam vad gäller dig."
"##emperor_favour_10##":"Kejsaren är fundersam vad gäller dig."
"##emperor_favour_11##":"Kejsaren tror du kan bevisa dig värdefull ."
"##emperor_favour_12##":"Kejsaren är tillfreds med dig."
"##emperor_favour_13##":"Kejsaren är mycket nöjd med vad du gjort."
"##emperor_favour_14##":"Kejsaren är mycket entusiastisk över vad du gjort."
"##emperor_favour_15##":"Kejsaren är nöjd med vad du gjort."
"##emperor_favour_16##":"Kejsaren är entusiastisk över vad du gjort."
"##emperor_favour_17##":"Kejsaren är extremt entusiastisk över vad du gjort."
"##emperor_favour_18##":"Kejsaren är utom sig av glädje över vad du gjort."
"##emperor_favour_19##":"Kejsaren är mer än tillfreds med vad du gjort."
"##emperor_favour_20##":"Kejsaren är så otroligt nöjd att han talar om att utnämna dig till sin arvinge."
"##emperor_request##":"Kejserlig begäran"
"##emperor_send_money_to_you_nearest_time##":"Det faktum att kejsaren nyligen måste ingripa för att rädda dig skadar allvarligt din stads rykte om välstånd."
"##emperor_wrath_by_debt_text##":"Jag är mycket missnöjd. Trots alla pengar jag har investerat i din stad och senatens generösa krediter, har du svikit mig. Din stad har inte betalat tillbaka sina lån. Mitt förtroende för dig var missriktat och jag tvingas nu finna en annan ståthållare i ditt ställe. Du kanske passar bättre i den nya position jag har i åtanke för dig..."
"##emperor##":"Imperiet"
"##emperoradv_caesar_has_high_respect_for_you##":"Caesar respekterar dig mer än någon annan ståthållare någonsin!"
"##emperror_legion_at_out_gates##":"En legion av kejsarens trupper står vid portarna"
"##empire_map##":"Gå till imperiet"
"##empire_service_tip##":"Sänd iväg trupper för att skydda"
"##empire_tax##":"Tribut"
"##empireBtnTooltip##":""
"##empiremap_our_city##":"Vår stad!"
"##employee##":"Enhet"
"##employees##":"Enheter"
"##employers##":"Anställd arbetsstyrka"
"##empmap_distant_romecity_tip##":"Avlägsen romersk stad"
"##emw_bought##":"Köpt"
"##emw_buy##":"Inköp"
"##emw_sell##":"Försäljningar"
"##emw_sold##":"Sålt"
"##enemy_army_threating_a_city##":"En fiendearmé som hotar en av rikets städer"
"##engineer_average_life##":"Allt tycks fungera väl här."
"##engineer_building_allok##":"Jag behövs knappast. Dessa byggnader är i utmärkt skick."
"##engineer_gods_angry##":"Måtte gudarna vara mig nådiga. Det är inte mitt fel att ståthållaren hånar dem."
"##engineer_good_life##":"Var hälsad! Är det inte en fantastisk stad?"
"##engineer_have_trouble_buildings##":"Dessa byggnader är i dåligt skick. Jag kom precis i rätt tid."
"##engineer_high_workless##":"Jag har tur som har ett arbete i denna tid av arbetslöshet."
"##engineer_low_entertainment##":"Efter en hård dags arbete vill jag se en bra pjäs eller strid. Det finns inte mycket chans till det i den här staden."
"##engineer_need_workers##":"Staden skulle fungera bättre om det fanns nog med arbetare."
"##engineer_salary##":"Ingenjörslön på"
"##engineer_so_hungry##":"Om jag inte får mat snart ger jag mig av från staden."
"##engineer##":"Ingenjör"
"##engineerBtnTooltip##":""
"##engineering_post_bad_work##":"Vi arbetar med minimistyrka. Vi kan knappt sända ut en ingenjör per månad på fältet."
"##engineering_post_full_work##":"För närvarande har vi inga driftavbrott Våra ingenjörer är alltid ute och inspekterar och reparerar skador på stadens byggnader."
"##engineering_post_info##":"Ingenjörer är mycket respekterade yrkesmän, och det är alltid stor efterfrågan på deras tjänster. Konstant underhåll förhindrar att byggnaderna faller samman."
"##engineering_post_need_some_workers##":"Det tar en eller två dagar innan våra utarbetade ingenjörer är tillbaka på gatorna."
"##engineering_post_no_workers##":"Vi har inga ingenjörer anställda, och vår egen kontorsbyggnad riskerar att falla samman."
"##engineering_post_on_patrol##":"Vår ingenjör är ute och arbetar."
"##engineering_post_patrly_workers##":"Vi har för lite personal, så vi måste vänta en vecka innan våra ingenjörer är tillbaka i tjänst."
"##engineering_post_ready_for_work##":"Vår ingenjör förbereder sig för att ge sig av."
"##engineering_post_slow_work##":"Vi är kraftigt underbemannade och har en tidslucka på två veckor mellan ingenjörernas rundor."
"##engineering_post##":"Ingenjörspostering"
"##engineering_structures##":"Ingenjörsbyggnader"
"##entadv_small_city_not_need_entert##":"För tillfället har dina medborgare enklare bestyr än underhållning att tänka på. Men i takt med att staden växer kommer de att begära något som lindrar monotonin i deras vardagsliv."
"##enter_your_name##":"Välj ett namn"
"##entertainment_advisor_title##":"Underhållning"
"##entertainment_need_for_upgrade##":"I delar av staden klagar man över frånvaron av fritidsanläggningar. Byggnation av fler platser för underhållning skulle hjälpa utvecklingen i de fattigare områdena."
"##entertainment_short##":"Ent"
"##entertainment##":"Underhållning"
"##entertainmentBtnTooltip##":""
"##etertadv_as_city_grow_you_need_more_entert##":"Medborgare som söker tidsfördriv har allt vad de behöver. Men i takt med att staden växer måste du förse dem med mer storslagen form av underhållning."
"##exit_point##":"Utträdespunkt"
"##exit_salary_window##":"Lämna löneskärmen"
"##exit_this_panel##":"Avsluta denna panel"
"##exit_without_saving_question##":"Var försiktig med att riva broar. Isolerade samhällen går snabbt under om de skärs av från vägen till Rom."
"##exit##":"Avsluta"
"##explosion##":"Explosion"
"##export_btn_tooltip##":"Fastställ den kvantitet av dessa varor som du önskar behålla innan de exporteras"
"##exports_over##":"Exportera vara över"
"##extreme_fire_risk##":"Extrem brandrisk"
"##factory_need_more_workers##":"Fungerar knappt. Tilldela fler människor till vår sektor"
"##farm_need_farmland##":"Bygg jordbruk på jordbruksmark (leta efter gult gräs)"
"##farm_working_bad##":""
"##farm_working_normally##":""
"##farm##":"Lantbruk"
"##favor_rating##":"Popularitetsställning"
"##favor##":"Popularitet"
"##festivals##":"Festivaler"
"##few_crime_risk##":"Detta är ett område med låg brottslighet, men vissa boende har klagat"
"##fig_farm_bad_work##":"Mycket få människor arbetar i denna fruktträdgård. Fruktskörden kommer att bli liten och sen."
"##fig_farm_full_work##":"Denna fruktträdgård har alla anställda den behöver. Träden dignar av mogen frukt."
"##fig_farm_info##":"Frukt är en viktig del av den balanserad diet som ditt folk behöver för hälsa och glädje. I sädesmagasinen lagras frukt för lokal konsumtion, och i handelsmagasinen förvaras överskottet för export."
"##fig_farm_need_some_workers##":"Denna fruktträdgård är underbemannad. Den producerar mindre frukt än vad den borde."
"##fig_farm_no_workers##":"Denna fruktträdgård har inga anställda. Produktionen har upphört."
"##fig_farm_patrly_workers##":"Denna fruktträdgård utnyttjar inte maximal kapacitet. Som resultat kommer fruktproduktionen att gå långsammare."
"##fig_farm##":"Fruktodling"
"##file##":"Arkiv"
"##fileload_load_tlp##":"Öppna detta sparade spel"
"##finance_advisor##":"Stadens kapital"
"##finance_advisor##":"Finanser"
"##finances##":"Finanser"
"##fire##":"Brand"
"##fired##":"Avskedad!"
"##fishing_boat##":"Fiskebåt"
"##fishing_waters##":""
"##fishing_wharf##":"Fiskehamn"
"##floatsam_enabled##":"Vrakgods på?"
"##floatsam##":"Vrakgods"
"##for_second_year_broke_tribute##":"För andra året i rad har du inte betalat tribut till Rom. Detta håller på att bli ett stort problem för din framtida karriär."
"##fort_has_been_cursed_by_mars##":"Detta fort har förbannats av Mars. Det kommer att dröja innan några soldater vågar sig tillbaka hit."
"##fort_horse##":"Stödtrupp - Ridande"
"##fort_info##":"Ett romerskt fort rekryterar soldater från förläggningar. Lägga till en militärhögskola skulle ge trupper med bättre utbildning."
"##fort_javelin##":"Kastspjut"
"##fort_legionaries_no_workers##":"Utan personal kan vi inte utbilda en enda ny rekryt. Mars hjälpe oss i krigstid!"
"##fort_legionaries##":"Legionärfort"
"##fort##":"Fort"
"##fortification_info##":"Murar saktar ner fiendens framstöt mot en stad. Murar kan raseras. Tjockare murar är starkare och dessutom ges vaktposterna i anslutna torn möjlighet att patrullera dem."
"##fortification##":""
"##forum_1_on_patrol##":"Vår indrivare är ute på inspektion."
"##forum_1_ready_for_work##":"Vår indrivare förbereder sig för att ge sig av."
"##forum_1_slow_work##":"Vi är kraftigt underbemannade och har en lucka på två veckor innan indrivarna ger sig ut."
"##forum_full_work##":"För närvarande arbetar våra indrivare med maximal effektivitet, och de är alltid ute och kontrollerar att alla förfallna skatter betalas in till staden."
"##forum_information##":"En populär samlingsplats och eftertraktat samhällselement. Forum anställer även skatteindrivare och är livsviktiga för stadens skattkammare."
"##forum_need_some_workers##":"Vi har korta avbrott i verksamheten, ungefär en dag eller två, innan våra indrivare är tillbaka på gatorna igen."
"##forum_no_workers##":"Utan indrivare bidrar det här kontoret inte med någonting till stadskassan."
"##forum_patrly_workers##":"Vi är underbemannade och måste vänta en vecka innan våra indrivare är tillbaka i tjänst."
"##forum##":"Forum"
"##fountain_info##":"Människorna hämtar allt vatten som de behöver från fontäner, som måste förses med vatten via ledningar från en reservoar. Fontäner är den källa till vatten som folket föredrar."
"##fountain_not_work##":"Denna fontän fungerar inte eftersom det inte finns tillräckligt med arbetare för att driva den."
"##fountain_will_soon_be_hooked##":"Denna fontän väntar på att anslutas till det underjordiska rörledningsnätet."
"##fountain##":"Fontän"
"##free##":"ledig"
"##freehouse_caption##":"Ledig tomt"
"##freehouse_text_noroad##":"Ingen kommer att skapa sig ett hem här eftersom det ligger för långt från närmaste väg. Om ingen väg byggs snart kommer detta område att återgå till öppet landskap."
"##freehouse_text##":"Ingen har så mycket som satt upp ett tält här ännu, fast immigranter kommer säkert att anlända inom kort om staden har tillgång till livsmedel och arbetstillfällen."
"##freespace_for##":"Utrymme för"
"##fruit_farm_slow_work##":"Med få anställda vid denna fruktträdgård kommer den lilla mängd frukt som mognar att ruttna bort."
"##fruit##":"Frukt"
"##fullscreen_off##":"Fönsterskärm"
"##fullscreen_on##":"Fullskärm"
"##funds_tooltip##":""
"##furniture_need##":"Möbler behövs"
"##furniture_workshop_bad_work##":"Med så få yrkesmän i snickeriet står produktionen nästan stilla. Det kommer inte att produceras mycket möbler under det kommande året."
"##furniture_workshop_full_work##":"Detta snickeri har full sysselsättning, och arbetar fullt ut med att producera möbler."
"##furniture_workshop_info##":"Snickarna vid snickeriet skapar fina möbler av virke. Medborgarna kan möblera sina villor och du kan handla med överskottet."
"##furniture_workshop_need_resource##":"Detta snickeri behöver leverans av virke från ett magasin eller från en brädgård för att kunna producera möbler."
"##furniture_workshop_need_some_workers##":"Detta snickeri är underbemannat, och det tar längre tid att producera möbler än vad det borde."
"##furniture_workshop_no_workers##":"Denna smedja har inga anställda. Produktionen har upphört."
"##furniture_workshop_patrly_workers##":"Detta snickeri har lediga platser. Möbelproduktionen blir snabbare när de besätts."
"##furniture_workshop_slow_work##":"Mycket få snickare arbetar här. Som resultat är möbelproduktionen långsam."
"##furniture_workshop##":"Möbelsnickeri"
"##furniture##":"Möbler"
"##game_is_paused##":"Spelet stoppat (Tryck P för att fortsätta)"
"##game_sound_options##":""
"##game_speed_options##":""
"##garden_info##":"Denna trevliga plats skänker medborgarna avkoppling från stadens buller, värme och smuts genom en sval oas av grönska. Alla vill ha en trädgård intill sitt hus."
"##garden##":"Trädgårdar"
"##gardens_info##":"Trädgårdar förbättrar den lokala miljön."
"##gatehouse##":"Grindstuga"
"##getting_reports_about_enemies##":"Vi får rapporter om fiender som närmar sig staden"
"##give_money_tip##":"Klicka här för att donera pengar till staden"
"##give_money##":"Ge pengar"
"##gladiator_gods_angry##":"Var hälsad, medborgare. Har du hört? Gudarna är vreda."
"##gladiator_good_life##":"Var hälsad. Livet här är skönt att leva, inte sant?"
"##gladiator_high_workless##":"De arbetslösa är så många här. Jag önskar vi kunde få träna oss på några av dem."
"##gladiator_low_entertainment##":"Tråkigt! Det säger alla om det här stället, trots mina tappra insatser. Staden behöver verkligen mer underhållning."
"##gladiator_need_workers##":"Det är hemskt. Jag har aldrig sett så många lediga jobb."
"##gladiator_perfect_life##":"Medborgare! Jag har kämpat i många städer och den här är en av de bästa."
"##gladiator_pit_bad_work##":"Jag har ingen personal utöver mig själv. Jag kan inte arbeta under dessa förhållanden! Som bäst kan jag utbilda en gladiator var tredje månad."
"##gladiator_pit_full_work##":"Det är med nöje vi tillkännager att vi, med full sysselsättning, utbildar upp till fyra nya gladiatorer varje månad."
"##gladiator_pit_need_some_workers##":"Vi är något underbemannade, och kan därför endast utbilda två nya gladiatorer i månaden."
"##gladiator_pit_no_workers##":"Utan utbildningspersonal kan denna skola inte utbilda nya gladiatorer."
"##gladiator_pit_patrly_workers##":"Vi har bara halva personalstyrkan, och kan därför endast utbilda en gladiator under nästa månad."
"##gladiator_pit_slow_work##":"Vi lider av svår personalbrist, och kommer att få kämpa för att utbilda en ny gladiator under de kommande två månaderna."
"##gladiator_pit##":"Gladiatorskola"
"##gladiator_so_hungry##":"Jag är så hungrig att jag kan äta ett lejon!"
"##gmenu_about##":"Om"
"##gmenu_advisors##":""
"##gmenu_exit_game##":"Avsluta spel"
"##gmenu_file_exit##":""
"##gmenu_file_mainmenu##":""
"##gmenu_file_restart##":""
"##gmenu_file_save##":""
"##gmenu_file##":""
"##gmenu_help##":""
"##gmenu_options##":""
"##gmsndwnd_ambient_sound##":"Ljudeffekter"
"##gmsndwnd_game_volume##":"Volym"
"##gmsndwnd_theme_sound##":"Musiken"
"##gmspdwnd_autosave_interval##":"Spara automatiskt varje månad"
"##gmspdwnd_game_speed##":""
"##gmspdwnd_scroll_speed##":""
"##go_to_problem##":"Klicka här för att gå till detta problemområde"
"##go2_problem_area##":"Gå till problemområde."
"##god_ceres_short##":"Ceres"
"##god_charmed##":"Charmerade"
"##god_displeased##":"Missnöjda"
"##god_exalted##":"Begeistrade"
"##god_excellent##":"Utmärkt"
"##god_good##":"Bra"
"##god_happy##":"Glada"
"##god_indifferent##":"Likgiltiga"
"##god_irriated##":"Sårade"
"##god_mars_short##":"Mars"
"##god_mercury_short##":""
"##god_neptune_short##":""
"##god_pleased##":"Nöjda"
"##god_poor##":"Dålig"
"##god_quitepoor##":"Mycket dålig"
"##god_veryangry##":"Vredgade"
"##god_verygood##":"Mycket bra"
"##god_verypoor##":"Mycket dålig"
"##god_wrathful##":"Rasande"
"##goth_warrior##":"En gotisk soldat"
"##goto_empire_map##":"Gå till kartan över imperiet"
"##goto##":"Gå till"
"##governor_palace_1_info##":"Ditt hem är en av stadens mest åtråvärda adresser. Dess storlek avgör hur stort välstånd vår stad kan uppnå."
"##governor_palace_1##":"Ståthållarens hus"
"##governor_palace_2##":"Ståthållarens villa"
"##governor_palace_3##":"Ståthållarens palats"
"##governor_salary_title##":"Personlig inkomst"
"##granaries_holds##":"månader"
"##granary_devastation_mode_text##":"Försöker att sända mat till annan plats"
"##granary_holds##":"månad"
"##granary_info##":"Fulla sädesmagasin är livsviktiga för att hålla folkets magar fyllda och för att attrahera nya medborgare. Ett sädesmagasin kan lagra säd, kött, grönsaker och frukt."
"##granary_orders##":"Instruktioner sädesmagasin"
"##granery##":"Sädesmagasin"
"##grape_factory_stock##":"Lagrade druvor,"
"##grape##":"Vindruvor"
"##graphics##":""
"##grass##":"Gräs"
"##great_festival##":"Storslagen festival"
"##greatPalace_info##":"De boende i detta palats befinner sig högst upp i det romerska samhället. De saknar inte något. Bara att lyckas hålla dem nöjda är en storartad insats."
"##greek_soldier##":"En grekisk soldat"
"##have_food_for##":"Livsmedelsförråd för"
"##have_less_academy_in_city_0##":"Du har för få högskolor i din stad. Om du bygger fler förbättras din ställning."
"##have_less_library_in_city_0##":"Du har för få bibliotek i din stad. Om du bygger fler förbättras din ställning."
"##have_less_school_in_city_0##":"Du har för få skolor i din stad. Om du bygger fler förbättras din ställning."
"##have_less_temple_in_city_0##":"Du har för få religiösa byggnader i din stad. Om du bygger fler förbättras din ställning."
"##have_less_theater_in_city_0##":"Du har för få teatrar i din stad. Om du bygger fler förbättras din ställning."
"##have_no_access_school_colege##":"Vissa områden kräver bättre tillgång till skolor och högskolor. Endast vissa hus har tillgång till skolor eller högskolor, och detta hindrar områdenas utveckling."
"##have_no_access_to_library##":"Tillgång till bibliotek krävs nu i vissa delar av staden. Dina medborgare har tid att läsa. Nu behöver de tillgång till litteratur."
"##have_no_food_on_next_month##":"- inga livsmedel kommande månad"
"##have_no_legions##":"Du har inga legioner att sända"
"##have_no_requests##":"För närvarande har du inga meddelanden att läsa. I takt med att din stad växer, eller om kejsaren begär varor av dig, kommer meddelanden att visas här"
"##having_some_slums_lack_migration##":"Att ha slumområden förhindrar immigration"
"##health_advisor##":"Hälsosituation"
"##health_advisor##":"Byggnader förknippade med hälsa"
"##health##":"Hälsa"
"##healthadv_noproblem_small_city##":"Din lilla bosättning har ännu inga hälsoproblem att rapportera."
"##healthadv_not_need_health_service_now##":"För närvarande finns ingen efterfrågan på hälsovård eller sanitära inrättningar. I takt med att staden utvecklas kommer dock befolkningen att kräva badhus och sjukhus, och senare även barberare!"
"##healthadv_some_regions_need_barbers_2##":"Vissa välbeställda delar av staden vill ha barberare. En lokal barberare ger bättre status åt området."
"##healthadv_some_regions_need_barbers##":"Fler områden i staden kräver nu barberare. I takt med att din stad blir allt mer välbeställd kommer fler att ha tid till rakning och klippning!"
"##healthadv_some_regions_need_bath_2##":"Vissa områden i staden behöver nu tillgång till badhus. Bristen på dessa sanitära anläggningar begränsar byggnadstillväxten i dessa områden."
"##healthadv_some_regions_need_bath##":"Vissa delar av staden vill ha fler badhus. Vissa hus har tillgång till bad, men andra har det inte, och detta hindrar deras utveckling."
"##healthadv_some_regions_need_doctors_2##":"Fler och fler människor vill ha bekväm tillgång till hälsovård. Anordna lokal tillgång till kliniker så att staden kan växa."
"##healthadv_some_regions_need_doctors##":"Vissa delar av staden kräver tillgång till en klinik. Utan någon form av hälsovård kommer dessa hus förmodligen inte att växa."
"##healthadv_some_regions_need_hospital##":"Utvecklingen i vissa områden hålls tillbaka av för få sjukhus i staden. Nya sjukhus attraherar fler patricierklasser till staden."
"##healthBtnTooltip##":""
"##help##":"Hjälp"
"##hide_bigpanel##":"Göm sidopanelen, och utöka spelvyn"
"##high_bridge##":"Fartygsbro"
"##high_crime_risk##":"Detta område står i begrepp att explodera i upplopp."
"##high_crime_risk##":"Hela detta område är som en jäsande krutdurk! Brottsligheten är epidemisk, och uppror sannolika"
"##high_damage_risk##":"Stor risk att kollapsa"
"##high_fire_risk##":"Stor brandrisk"
"##high_salary_angers_senate##":"Den löjligt höga lön du betalar till dig själv upprör senaten. Hela Rom talar om din öppna girighet."
"##hippodrome_full_access##":"Detta hus har tillgång till hippodrom"
"##hippodrome_haveno_races##":"Inga kapplöpningar för närvarande"
"##hippodrome_no_access##":"Detta hus har inte tillgång till hippodromen"
"##hippodrome_no_workers##":"Inget rör sig i hippodromen. Utan arbetare ger den ingen underhållning åt lokalsamhället."
"##hippodrome##":"Hippodrom"
"##hippodromes##":"Hippodromer"
"##hold_ceres_festival##":"Anordna festival för Ceres"
"##hold_mars_festival##":"Anordna festival för Mars"
"##hold_mercury_festival##":"Anordna festival för Merkurius"
"##hold_neptune_festival##":"Anordna festival för Neptunus"
"##hold_venus_festival##":"Anordna festival för Venus"
"##hospital_full_access##":"Detta hus har tillgång till sjukhus"
"##hospital_full_work##":"Detta sjukhus används, och betjänar lokalsamhället."
"##hospital_info##":"Även om ingen vill bo i närheten av dem, räddar sjukhus liv. Staden borde ha tillräckligt med sängplatser för alla sina invånare."
"##hospital_no_access##":"Detta hus har inte tillgång till ett sjukhus"
"##hospital_no_workers##":"Detta sjukhus används inte, och är därför värdelöst för lokalsamhället."
"##hospital##":"Sjukhus"
"##hospitals##":"Sjukhus"
"##house_evolves_at##":"Denna boning kommer snart att utvecklas och få bättre status, som ett resultat av de förbättrade lokala villkoren."
"##house_food_only_for_month##":"Detta hus har matförråd som åtminstone kommer att räcka under den kommande månaden"
"##house_have_not_food##":"Detta hus har inget livsmedelsförråd"
"##house_have_some_food##":"Detta hus kommer snart att äta sig igenom sitt begränsade livsmedelsförråd"
"##house_no_troubles_with_food##":"Detta hus har inget problem med att skaffa den mat som krävs för att överleva"
"##house_not_registered_for_taxes##":"Detta hus befinner sig i en region utan skatteadministration, och betalar därför ingen skatt"
"##house_not_report_about_crimes##":"De boende har inte rapporterat någon brottslighet."
"##house_provide_food_themselves##":"Tältboende hämtar sin egen mat från omgivande marker."
"##houseBtnTooltip##":""
"##how_to_grow_prosperity##":"Ställningen har inte förändrats detta året. Att visa vinst i stadens årliga räkenskaper är det bästa sättet att förbättra välståndsställningen."
"##hun_warrior##":"En hunnersoldat"
"##immigrant_much_food_here##":"De påstår att det finns mat här. Är det en bra plats att bo på?"
"##immigrant_so_hungry##":"Om jag stannar längre dör jag. Det finns ingen mat någonstans."
"##immigrant_want_to_be_liontamer##":"Jag har hört att det finns arbete här. Jag vill bli lejontämjare."
"##immigrant_where_my_home##":"Jag är ny i staden. Vet du var man kan få tag i en bostad?"
"##imperial_request_cance_badly_affected##":"Den kejserliga begäran som du nyligen upphävde har skadat din ställning i Rom."
"##import_fn##":"Importer"
"##import##":"Importerar"
"##industry_disabled##":"Industri är AV"
"##industry_enabled##":"Industri är PÅ"
"##infobox_construction_comma_tip##":"TIPS: Använd komma och punkt för snabbflyttning genom dessa och andra objekt."
"##infobox_tooltip_exit##":""
"##infobox_tooltip_help##":""
"##initialize_animations##":""
"##initialize_constructions##":""
"##initialize_house_specification##":""
"##initialize_names##":""
"##initialize_religion##":""
"##initialize_walkers##":""
"##inland_lake_text##":"Denna insjö saknar kontakt med havet"
"##iron_factory_stock##":"Lagrat järn,"
"##iron_mine_bad_work##":"Med så få anställda står produktion nästan stilla. Det kommer att produceras mycket lite järn under det närmaste året."
"##iron_mine_collapse##":"Malmbrott kollapsar"
"##iron_mine_full_work##":"Detta brott har alla anställda det behöver, och arbetar fullt ut med att producera järn."
"##iron_mine_info##":"Bryt järn för att handla med, eller för att leverera till vapensmedjorna. Utrusta din armé med hemgjorda vapen, eller exportera dem till andra provinser."
"##iron_mine_need_some_workers##":"Detta brott utnyttjar inte maximal kapacitet. Malmbrytningen skulle vara mycket effektivare med fler arbetare."
"##iron_mine_no_workers##":"Detta brott har inga anställda. Produktionen har upphört."
"##iron_mine_patrly_workers##":"Detta brott är underbemannat. Det tar längre tid än normalt att producera järnet."
"##iron_mine_slow_work##":"Mycket få människor arbetar vid det här brottet. Som resultat är järnproduktionen långsam."
"##iron_mine##":"Malmbrott"
"##iron##":"Järn"
"##its_very_peacefull_province##":"Imperiet har aldrig förut skådat en stad med sådant lugn!"
"##judaean_warrior##":"En judéisk soldat"
"##labor##":"Arbetskraft"
"##landmerchant_good_deals##":"Jag älskar att komma hit. Affärerna går mycket bra."
"##landmerchant_noany_trade##":"Jag vet inte varför jag tar den här handelsvägen. De köper ingenting och de har inget de vill sälja till mig."
"##landmerchant_say_about_store_goods##":"Försiktigt! Jag önskar att arbetarna skulle ta det lugnt när de lastar mina djur med de varor jag nyss har köpt."
"##landmerchart_noany_trade2##":"Inget att byteshandla med här, passerar bara"
"##large_temple##":"Stort tempel"
"##large_temples##":"Stora tempel"
"##large##":"Stort"
"##last_year##":"Förra året"
"##lawless_area##":"Ett laglöst område. Människorna är vettskrämda."
"##layer_crime##":"Brott"
"##leave_empire?##":"Lämna det Romerska Riket?"
"##left_click_open_right_erase##":"Vänsterklicka på ett meddelande för att läsa. Högerklicka för att radera."
"##legion_formation_tooltip##":"Klicka här för att ändra legionens formation"
"##legion_haveho_soldiers_and_barracks##":"Denna legion har för närvarande inga soldater. Den existerar bara till namnet och utan förläggningar i staden kan den inte ta emot några nya trupper."
"##legion_haveho_soldiers##":"Denna legion har för närvarande inga soldater. Den existerar bara till namnet. Endast när nyligen utbildade trupper anländer från förläggningarna kommer den att förvandlas till en stridande enhet."
"##legion##":"Militär"
"##legionadv_no_legions##":"Du har inga legioner att leda. Du måste först bygga ett fort"
"##legionary_average_life##":"Jag slåss intill döden! Staden är trygg så länge jag lever!"
"##legionary_low_salary##":"Jag får inte tillräckligt bra betalt för att slåss!"
"##legions##":"Legioner"
"##lgn_heroes##":"Hjältarna"
"##lgn_hydras##":"Hydrorna"
"##lgn_lions##":"Lejonen."
"##lgn_pigs##":"Svinen"
"##lgn_rabbits##":"Kaninerna"
"##lgn_snakes##":"Ormarna"
"##lgn_stallion##":"Hingstarna"
"##lgn_wolves##":"Vargarna"
"##libraries##":"Bibliotek"
"##library_access_perfectrly##":"Områden som kräver utbildningsmöjligheter har tillgång till dem, men fler bibliotek skulle minska trängseln."
"##library_full_access##":"Detta hus har tillgång till bibliotek"
"##library_full_work##":"Detta bibliotek används. Dess hyllor är fyllda med skriftrullar med lärdom."
"##library_info##":"Litterära arbeten från hela riket förvaras här på grekiska och latin. Lärda män insisterar att biblioteken är avgörande för en viktig stad."
"##library_no_access##":"Detta hus har inte tillgång till bibliotek"
"##library_no_workers##":"Hyllorna i detta bibliotek är tomma, och värdelösa för lokalsamhället."
"##library##":"Bibliotek"
"##lindum_extremely_dangerous_province##":"Lindum: en extremt farlig provins"
"##lion_pit_bad_work##":"Jag har ingen personal utöver mig själv. Jag kan inte arbeta under dessa förhållanden! Som bäst kan jag leverera ett lejon på tre månader."
"##lion_pit_need_some_workers##":"Vi är något underbemannade, och kan därför endast leverera två nya lejon i månaden."
"##lion_pit_no_workers##":"Utan personal kan detta lejonhus inte leverera några nya lejon till spelen."
"##lion_pit_patrly_workers##":"Vi har bara halva personalstyrkan, och kan därför endast leverera ett lejon under nästa månad."
"##lion_pit_slow_work##":"Vi lider av svår personalbrist, och kommer att få kämpa för att leverera ett enda lejon under de kommande två månaderna."
"##lion_pit_work##":"Det är med nöje vi tillkännager att vi, med full sysselsättning, kan leverera upp till fyra nya lejon varje månad."
"##lion_pit##":"Lejonhus"
"##lionTamer_average_life##":"Här är lite utländskt kött åt dig, Leo."
"##lionTamer_gods_angry##":"Gudarna är så vreda att det påverkar mitt lejon. Han är vrålarg."
"##lionTamer_good_education##":"Var hälsad. Den här staden tycker vi om, inte sant, Leo?"
"##lionTamer_good_life##":"Nu har du din chans, Leo. Duktigt lejon."
"##lionTamer_high_workless##":"Det är stor arbetslöshet här."
"##lionTamer_low_entertainment##":"Leo och jag slåss dygnet runt och ändå har folk tråkigt. Det finns helt enkelt inte tillräckligt med artister här."
"##lionTamer_need_workers##":"Den här staden behöver mer arbetskraft. Jag undrar om jag kan träna Leo att arbeta mer?"
"##lionTamer_so_hungry##":"Om vi inte får mer mat snart, äter lejonet upp mig!"
"##little_damage_risk##":"Viss risk att kollapsa"
"##Load_save##":"Öppna sparat spel"
"##loading_offsets##":""
"##loading_resources##":" "
"##londinium_win_text##":"Vid Jupiter! Vildarna i Britannia har aldrig sett Londiniums like. Claudius, som visade öborna de romerska svärdens vassa eggar för många år sedan, ler säkert mot oss från sin himmel."
"##lost_money_last_year##":"Förra året förlorade din stad pengar - detta minskade stadens välstånd."
"##low_bridge##":"Låg bro"
"##low_crime_risk##":"Brott inträffar sällan i detta område"
"##low_damage_risk##":"Liten risk att kollapsa"
"##low_desirability_degrade##":"Detta hus kommer snart att förfalla. Den sjunkande efterfrågan på boende i detta område drar ner det."
"##low_desirability##":"Du behöver göra området mer attraktivt, t ex genom att anlägga några trädgårdar eller torg."
"##low_fire_risk##":"Liten brandrisk"
"##low_wage_broke_migration##":"Låga löner förhindrar immigration"
"##low_wage_broke_migration##":"Låga löner minskar immigrationen till din stad"
"##low_wage_lack_migration##":"Låga löner är ett problem"
"##lugdunum_win_text##":"Din behandling av gallerna i Lugdunum och den sköna stadens prakt bådar väl för Roms expansion i den norra vildmarken. Bra gjort!"
"##lumber_mill_bad_work##":"Det finns nästan inga skogsarbetare, och produktionen står nästan still."
"##lumber_mill_full_work##":"Denna brädgård har alla anställda den behöver. Den arbetar fullt ut med att såga timmer."
"##lumber_mill_info##":"Såga virke för handel, eller till möbelverkstäderna. Patricierna vill ha möbler till sina villor, eller så kan du exportera det till dina handelspartners."
"##lumber_mill_need_some_workers##":"Denna brädgård är underbemannad, och det tar längre tid att såga virke än vad det borde."
"##lumber_mill_need_some_workers##":"Denna brädgård arbetar inte med maximal kapacitet. Som resultat kommer timmerproduktionen att bli något långsammare."
"##lumber_mill_no_workers##":"Denna brädgård har inga anställda. Produktionen har upphört."
"##lumber_mill_slow_work##":"Mycket få människor arbetar vid den här brädgården. Som resultat är timmerproduktionen långsam."
"##lumber_mill##":"Brädgård"
"##lutetia_win_text##":"Kejsar Augustus måste ha anat ditt styre när han förutspådde vår seger över gallerna. Din framgång vid Lutetia räcker långt när det gäller att krossa deras upprorsanda."
"##luxury_palace##":"Lyxpalats"
"##macedonian_soldier##":"En makedonisk soldat"
"##mainmenu_credits##":"Credits"
"##mainmenu_language##":""
"##mainmenu_load##":"Öppna spel"
"##mainmenu_loadcampaign##":""
"##mainmenu_loadgame##":"Öppna spel"
"##mainmenu_loadmap##":"Ny karta"
"##mainmenu_newgame##":"Nytt spel"
"##mainmenu_options##":""
"##mainmenu_playmission##":""
"##mainmenu_quit##":"Avsluta spel"
"##mainmenu_randommap##":"Öppet spel "
"##mainmenu_sound##":"Ljud"
"##mainmenu_video##":"Bild"
"##marble##":"Marmor"
"##market_about##":"Våra marknader gör imperiets rika håvor tillgängliga för medborgare med pengar. Varje hem behöver tillgång till en marknad, men ingen vill bo intill en."
"##market_full_work##":"Denna marknad används"
"##market_kid_say_1##":"Den tjocka damen bad mig bära detta och följa efter henne."
"##market_no_workers##":"Denna marknad används inte, och levererar inga produkter till lokalsamhället."
"##market_search_food_source##":"Denna marknad har köpmän men de söker för närvarande efter en källa till livsmedel som kan säljas."
"##market##":"Marknad"
"##marketBuyer_average_life##":"Denna stad är egentligen inte så illa."
"##marketBuyer_find_goods##":"Jag ska hämta nya varor."
"##marketBuyer_gods_angry##":"Detta är en hednisk plats. Ståthållaren har ingen respekt för gudarna."
"##marketBuyer_good_life##":"God dag, medborgare. Är det inte en härlig stad?"
"##marketBuyer_high_workless##":"Med denna höga arbetslöshet måste jag arbeta hårt för att behålla mitt jobb."
"##marketBuyer_low_entertainment##":"Detta måste vara den tråkigaste staden i imperiet."
"##marketBuyer_need_workers##":"Jag har aldrig sett så många byggnader som behöver fler arbetare."
"##marketBuyer_return##":"Dessa korgar är så tunga! Jag har med mig färska varor till min marknad."
"##marketBuyer_so_hungry##":"Det finns inte tillräckligt med livsmedel här. Hur ska jag kunna försörja mig?"
"##marketKid_say_2##":"Korgen tar kål på mig. Jag bryr mig inte om vem som behöver maten, det borde finnas en lag mot barnarbete."
"##marketKid_say_3##":"Var hälsad! Jag bär korgen med mat till kvinnans marknad. Jag hoppas jag får bra med dricks!"
"##marketLady_no_food_on_market##":"Marknaden har slut på livsmedel, så jag är på väg hem."
"##mars_desc##":"Krig"
"##mars_watches_over_soldiers##":"Mars vakar över soldater och belönar tapperhet i fält. Ingen man vågar kämpa utan Mars välsignelse."
"##massilia_preview_mission##":"Det enda vattnet finns i oasen. Detsamma gäller tyvärr för odlingsbar mark. Reservoarer och lantgårdar konkurrerar om samma utrymme. Använd det med förstånd."
"##max_available##":"Underhåller"
"##maximizeBtnTooltip##":""
"##may_collect_about##":"ger en avkastning på"
"##meadow_caption##":"Äng"
"##meat_farm_bad_work##":"Det finns knappt några anställda vid den här farmen, och dess djurstam är liten och sjuklig."
"##meat_farm_full_work##":"Denna farm har alla anställda den behöver, och dess djurstam är fet och stor."
"##meat_farm_info##":"Välmående medborgare njuter av olika sorters fläsk. Kött kan förvaras i sädesmagasin för lokal konsumtion eller i handelsmagasin för export."
"##meat_farm_need_some_workers##":"Denna farm är underbemannad. Svinen har små kullar, som växer långsamt."
"##meat_farm_no_workers##":"Denna farm har inga anställda, och alla djuren har flytt eller dött."
"##meat_farm_patrly_workers##":"Denna farm arbetar inte med maximal kapacitet. Som resultat kommer köttproduktionen att bli något mindre."
"##meat_farm_slow_work##":"Mycket få människor arbetar på den här farmen. Som resultat är köttproduktionen långsam."
"##meat_farm##":"Svinuppfödning"
"##meat##":"Kött"
"##mediolanum_win_text##":"Att Hannibal kunde korsa Alperna med sina elefanter var häpnadsväckande. Att Mediolanum skulle blomstra trots hans attacker är ett mirakel. Din framgång vände lyckan i det puniska kriget till Roms fördel. Hela Rom tackar dig."
"##mercury_desc##":"Handel"
"##mercury##":"Mercury"
"##message##":"Meddelande"
"##messageBtnTooltip##":"Meddelanden från dina skrivare"
"##messages##":"Meddelanden"
"##middle_festival##":"Stor festival"
"##middle_file_risk##":"Denna byggnad har en viss brandrisk"
"##middle_insula##":"Medelstor Insulae"
"##middle_palace##":"Medelstort palats"
"##middle_villa##":"Medelstor villa"
"##migration_broke_tax##":"Höga skatter gör att vissa människor undviker din stad"
"##migration_broke_workless##":"Hög arbetslöshet i din stad bromsar din välståndsställning."
"##migration_empty_granary##":"Brist på mat förhindrar immigration"
"##migration_lack_crime##":"Hög brottslighet skrämmer lokalbefolkningen."
"##migration_lack_empty_house##":"Brist på husrum begränsar immigrationen"
"##migration_lack_tax##":"Höga skatter är ett problem"
"##migration_lack_workless##":"Arbetslöshet minskar antalet immigranter"
"##migration_lessfood_granary##":"Brist på livsmedel i sädesmagasinen minskar immigrationen"
"##migration_low_food_stocks##":"Bristen på mat är ett problem"
"##migration_middle_lack_tax##":"Höga skatter förhindrar immigration"
"##migration_middle_lack_workless##":"Hög arbetslöshet är ett problem"
"##migration_middle_lack_workless##":"Brist på arbete förhindrar immigration"
"##migration_people_away##":"Brist på arbete driver bort människor"
"##migration_war_deterring##":"Krig avskräcker immigranter!!"
"##miletus_win_text##":"Precis som jag förväntade mig har exemplet Miletus redan inspirerat andra östliga städer att inleda förhandlingar om att ingå i imperiet. Din erfarenhet av fisket har blivit en läxa för alla mina ståthållare!"
"##military_academy_patrly_workers##":"När nya soldater har avslutat sin utbildning i förläggningen kommer de hit för att förbättra och finslipa sina färdigheter. Det går dock först när vi har fått tillräckligt med personal."
"##militaryAcademy_full_work##":"Vi förser nya rekryter från stadens förläggningar med den ytterligare utbildning de kräver för att fungera bra i en modern romersk armé."
"##militaryAcademy_no_workers##":"Utan personal kan vi inte finslipa kunskaperna för stadens nya soldater. De tvingas att gå direkt till sina fort och sedan hoppas på det bästa..."
"##militaryAcademy##":"Militärhögskola"
"##minimap_tooltip##":"Klicka på denna översiktskarta för att flytta till avlägsna delar av din stad"
"##minimizeBtnTooltip##":""
"##missing_barber_degrade##":"Detta hus kommer snart att förfalla, eftersom det har förlorat tillgången till barberare."
"##missing_barber##":"Detta hus kan inte utvecklas, eftersom det inte har någon lokal tillgång till en barberare."
"##missing_bath_degrade##":"Detta hus kommer snart att förfalla, eftersom det har förlorat tillgången till sitt badhus."
"##missing_bath##":"Detta hus kan inte utvecklas, eftersom det inte har tillgång till ett lokalt badhus."
"##missing_college_degrade##":"Detta hus kommer snart att förfalla. Dess tidigare utmärkta tillgång till utbildning har försämrats, eftersom det har förlorat tillgången till sin högskola."
"##missing_college##":"Detta hus kan inte utvecklas, eftersom dess redan utmärkta tillgång till utbildning måste förbättras genom tillgång till en högskola."
"##missing_doctor__degrade##":"Detta hus kommer snart att förfalla, eftersom dess möjligheter till hälsovård skurits ned. Det finns lokal tillgång till ett sjukhus men det är svårt att hitta en klinik."
"##missing_doctor_or_hospital_degrade##":"Detta hus kommer snart att förfalla, eftersom det nu har tvivelaktig hälsovård. Det saknas inte bara tillgång till en klinik, utan även tillgången till sjukhus är dålig."
"##missing_doctor_or_hospital##":"Detta hus kan inte utvecklas, eftersom det i stort sett saknar tillgång till sjukvård. Det saknar tillgång till både klinik och sjukhus."
"##missing_doctor##":"Detta hus kan inte utvecklas, eftersom det vill ha bättre möjligheter till sjukvård. Det finns lokal tillgång till ett sjukhus men det behövs en klinik i närheten."
"##missing_entertainment_also_degrade##":"Detta hus kommer snart att förfalla. Det finns god underhållning i området, men inte tillräckligt varierat utbud."
"##missing_entertainment_also##":"Detta hus kan inte utvecklas, eftersom det inte finns tillräckligt med underhållning i området."
"##missing_entertainment_amph_degrade##":"Detta hus kommer snart att förfalla. Det finns viss underhållning i området, men inte tillräckligt."
"##missing_entertainment_amph##":"Detta hus kan inte utvecklas, eftersom det knappt finns någon underhållning i området."
"##missing_entertainment_colloseum_degrade##":"Detta hus kommer snart att förfalla. Det finns utmärkt underhållning i området, men det är trångt och utbudet är inte tillräckligt varierat för de kräsna patricierna."
"##missing_entertainment_colloseum##":"Detta hus kan inte utvecklas, eftersom det visserligen finns viss underhållning i området, men inte tillräckligt."
"##missing_entertainment_degrade##":"Detta hus kommer snart att förfalla, eftersom det knappast finns någon underhållning i området."
"##missing_entertainment_degrade##":"Detta hus kommer snart att förfalla, eftersom det inte finns tillräckligt med underhållning i området."
"##missing_entertainment_need_more##":"Detta hus kan inte utvecklas, eftersom det visserligen finns god underhållning i området, men inte tillräckligt varierat utbud."
"##missing_entertainment_patrician##":"Detta hus kan inte utvecklas, eftersom det visserligen finns utmärkt underhållning i området, men det är trångt och utbudet är inte tillräckligt varierat för de kräsna patricierna."
"##missing_entertainment##":"Detta hus kan inte utvecklas, eftersom det inte finns någon underhållning i området."
"##missing_food_degrade##":"Detta hus kommer snart att förfalla, eftersom det inte har fått några livsmedelsleveranser från en lokal marknad nyligen."
"##missing_food_degrade##":"Detta hus kommer snart att förfalla. Det har visserligen tillgång till en marknad, men marknaden själv har svårt att få livsmedelsleveranser."
"##missing_food_from_market##":"Detta hus kan inte utvecklas. Det har visserligen tillgång till en lokal marknad, men marknaden själv har svårt att få livsmedelsleveranser."
"##missing_food##":"Detta hus kan inte utvecklas, eftersom det måste ha leveranser av livsmedel från en lokal marknad."
"##missing_fountain_degrade##":"Detta hus kommer snart att förfalla, eftersom det inte har tillgång till rent vatten från en fontän."
"##missing_fountain##":"Detta hus kan inte utvecklas, eftersom det inte har tillgång till ren vattentillförsel från en fontän."
"##missing_furniture_degrade##":"Detta hus kommer snart att förfalla, eftersom det har slut på möbler och dess lokala marknad har ett sporadiskt utbud."
"##missing_furniture##":"Detta hus kan inte utvecklas. Det behöver tillgång till möbelleveranser från sin lokala marknad innan mer välmående medborgarklasser kommer att flytta in."
"##missing_hospital_degrade##":"Detta hus kommer snart att förfalla, eftersom dess tillgång till hälsovård har skurits ned. Tillgången till kliniker är god men det finns inga lokala sjukhus."
"##missing_hospital##":"Detta hus kan inte utvecklas, eftersom det vill ha bättre möjligheter till sjukvård. Klinikernas täckning är bra men det saknas lokal tillgång till ett sjukhus."
"##missing_library_degrade##":"Detta hus kommer snart att förfalla. Dess tillgång till utbildning har försämrats, eftersom det har förlorat tillgång till sitt bibliotek."
"##missing_library##":"Detta hus kan inte utvecklas, eftersom dess tillgång till utbildning måste förbättras genom tillgång till ett bibliotek."
"##missing_market_degrade##":"Detta hus kommer snart att förfalla. Det har förlorat tillgången till en marknad."
"##missing_market##":"Detta hus kan inte utvecklas, eftersom det inte har tillgång till en lokal marknad."
"##missing_oil_degrade##":"Detta hus kommer snart att förfalla, eftersom det har slut på oljan och dess lokala marknad har ett sporadiskt utbud."
"##missing_oil##":"Detta hus kan inte utvecklas. Det behöver oljeleveranser från sin lokala marknad innan mer välmående medborgarklasser kommer att flytta in."
"##missing_pottery_degrade##":"Detta hus kommer snart att förfalla. Det har inte längre tillgång till krukor, och leveranserna till dess lokala marknad är minst sagt opålitliga."
"##missing_pottery##":"Detta hus kan inte utvecklas. Det behöver leveranser av krukor från sin lokala marknad innan förmögnare medborgarklasser kommer att flytta in."
"##missing_religion_degrade##":"Detta hus kommer snart att förfalla, eftersom det har förlorat all tillgång till lokala religiösa byggnader."
"##missing_religion##":"Detta hus kan inte utvecklas, eftersom det inte har tillgång till några lokala möjligheter till religionsutövning."
"##missing_school_degrade##":"Detta hus kommer snart att förfalla. Dess tillgång till utbildning har försämrats, eftersom det har förlorat tillgång till sin skola."
"##missing_school_or_library_degrade##":"Detta hus kommer snart att förfalla, eftersom det har förlorat alla grundläggande utbildningsmöjligheter från en skola eller ett bibliotek."
"##missing_school_or_library##":"Detta hus kan inte utvecklas, eftersom det inte har tillgång till grundläggande utbildningsmöjligheter vare sig från skola eller bibliotek."
"##missing_school##":"Detta hus kan inte utvecklas, eftersom dess tillgång till utbildning måste förbättras genom tillgång till en skola."
"##missing_second_food_degrade##":"Detta hus kommer snart att förfalla, eftersom det endast har tillgång till en enda typ av livsmedel från sin lokala marknad. Detta avskräcker de välbärgade klasserna."
"##missing_second_food##":"Detta hus kan inte utvecklas, eftersom det krävs en till typ av livsmedel, som levereras från en lokal marknad, för att förmå mer välbärgade att flytta in."
"##missing_second_religion_degrade##":"Detta hus kommer snart att förfalla. Dess tillgång till lokala religiösa byggnader har reducerats till endast ett tempel för en enda gud."
"##missing_second_religion##":"Detta hus kan inte utvecklas, eftersom det endast har tillgång till tempel för en enda gud. I takt med att dess invånare kommer upp sig i världen kommer de att vilja ägna mer tid åt att tillbe andra gudar."
"##missing_second_wine##":"Detta hus kan inte utvecklas. Det krävs en vinsort till för att tillfredsställa de sysslolösa patriciernas dekadenta livsstil. Öppna en ny handelsväg, eller tillverka ditt eget vin."
"##missing_third_food_degrade##":"Detta hus kommer snart att förfalla, eftersom det endast har tillgång till 2 typer av livsmedel från sin lokala marknad. Detta avskräcker patricierklasserna."
"##missing_third_food##":"Detta hus kan inte utvecklas, eftersom det krävs en tredje typ av livsmedel, som levereras från en lokal marknad, för att förmå patricierklasserna att flytta in."
"##missing_third_religion_degrade##":"Detta hus kommer snart att förfalla. Dess tidigare utmärkta religiösa möjligheter har reducerats, och det har nu endast tillgång till tempel för två gudar."
"##missing_third_religion##":"Detta hus kan inte utvecklas, eftersom det endast har tillgång till tempel för två gudar. I takt med att dess invånare kommer upp sig i världen kommer de att vilja ägna mer tid åt att tillbe andra gudar."
"##missing_water_degrade##":"Detta hus kommer snart att förfalla, eftersom det saknar tillgång till även den enklaste vattenförsörjning."
"##missing_water##":"Detta hus kan inte utvecklas, eftersom det inte har tillgång till ens den mest primitiva vattenförsörjning."
"##missing_wine_degrade##":"Detta hus kommer snart att förfalla, eftersom det har slut på vin och dess lokala marknad har ett sporadiskt utbud."
"##missing_wine##":"Detta hus kan inte utvecklas. Det behöver tillgång till vinleveranser från sin lokala marknad innan mer välmående medborgarklasser kommer att flytta in."
"##mission_win##":"Seger"
"##mission_wnd_population##":"Befolkning"
"##mission_wnd_targets_title##":"Mål"
"##mission_wnd_tocity##":"Till staden"
"##missionaryPost_full_work##":"Vi arbetar på att civilisera lokalbefolkningen. Genom att lära dem grunderna i latin hoppas vi uppmuntra dem att arbeta med oss, istället för emot oss."
"##missionaryPost##":"Inhemsk mission"
"##missionBtnTooltip##":"Titel på provinskarta."
"##moment_fire_risk##":"Denna byggnad kan fatta eld när som helst!"
"##month_1_short##":"Jan"
"##month_10_short##":"Okt"
"##month_11_short##":"Nov"
"##month_12_short##":""
"##month_2_short##":""
"##month_3_short##":"Mar"
"##month_4_short##":""
"##month_5_short##":"Maj"
"##month_6_short##":"Jun"
"##month_7_short##":"Jul"
"##month_8_short##":""
"##month_9_short##":"Sep"
"##month_from_last_festival##":"sedan senaste festivalen"
"##month##":"Person"
"##months_until_defeat##":"månader till nederlag"
"##months_until_victory##":"månader till seger"
"##months##":"Människor"
"##more_0_month_from_festival##":"Ditt folk, somliga fortfarande berusade efter festen, välkomnar din generositet."
"##more_12_month_from_festival##":"Ditt invånare är mycket missnöjda med tanken på ännu ett år utan en festival."
"##more_16_month_from_festival##":"Människorna kommer inte längre ihåg den sista festivalen som hölls i staden."
"##more_4_month_from_festival##":"Människor talar fortfarande varmt om din senaste festival."
"##more_8_month_from_festival## ":"Minnet av den tidigare festivalen håller på att blekna."
"##more_people##":"Anställda"
"##more_person##":"Anställd"
"##more_salary_dispeasure_senate##":"Den lön som du betalar dig själv, och som vida överskrider din rang, är en källa till missnöje i Rom."
"##much_plebs##":"Den höga koncentrationen av boende i slumområden i din stad gör att den ser fattig ut."
"##my_rome##":""
"##nativeCenter_info##":"Mötesplatsen för den lokalbefolkning som kommer hit för att byteshandla med enkla handelsvaror. Om styresmannen bara kunde lära sig några ord på latin..."
"##nativeCenter##":"Inhemskt centrum"
"##nativeField_info##":"Vissa primitiva grödor, som förser lokalbefolkningen med en grundläggande källa till livsmedel."
"##nativeField##":""
"##nativeHut_info##":"En del lokalbefolkning bor här, de lever ett stillsamt enkelt liv. De vill bara bli lämnade ifred."
"##nativeHut##":"Infödingshydda"
"##nearby_building_negative_effect_degrade##":"En närliggande byggnad har en försämrande effekt på efterfrågan till området. Försök att anlägga t ex trädgårdar, torg och statyer."
"##nearby_building_negative_effect##":"En närliggande byggnad har en försämrande effekt på efterfrågan till området. Försök att anlägga t ex trädgårdar, torg och statyer."
"##need_access_to_full_reservoir##":"Kräver tillgång till en full reservoar för att fungera"
"##need_actor_colony##":"Bygg en skådespelarkoloni för att sända skådespelare hit"
"##need_barracks_for_work##":"Fungerande förläggning krävs för att ta emot soldater"
"##need_build_on_cleared_area##":"Måste byggas på avröjt land"
"##need_build_on_cleared_area##":""
"##need_charioter_school##":"Bygg en skola för körsvenner för att se kapplöpningar"
"##need_clay_pit##":"Denna byggnad kräver lera"
"##need_grape##":"Denna byggnad kräver druvor"
"##need_iron_for_work##":"Denna byggnad kräver järnmalm"
"##need_iron_mine##":"Bygg en järngruva"
"##need_lionnursery##":"Bygg ett lejonhus för att arrangera djurtävlingar"
"##need_marble_for_large_temple##":"Du behöver 2 ton marmor för att bygga ett stort tempel"
"##need_olive_farm##":"Bygg en olivodling"
"##need_population##":"krävs)"
"##need_reservoir_for_work##":"Denna fontän fungerar inte eftersom den inte ligger i ett område som täcks av rörledningar från en fungerande reservoar."
"##need_temples_for_city##":"Dina medborgare har börjat bli intresserade av religion. Frånvaron av en närliggande gudstjänstplats hindrar stadens utveckling."
"##need_timber_mill##":"Bygg en brädgård"
"##need_trainee_charioteer##":"Det finns inga kapplöpningsvagnar i din hippodrom. Anskaffning av sådana skulle avsevärt förbättra villkoren för befolkningen, som ivrigt söker mer underhållning."
"##need_vines_farm##":"Bygg en vingård"
"##neptune_desc##":"Havet"
"##neptune_despleasure_tip##":"Sjömän finner att Neptunus är en ombytlig gud även om han blidkas. Väck inte Neptunus vrede, om du önskar bedriva handel över vattnet."
"##neptune_wrath_of_you##":"Neptunus skyddar sjömän och deras skepp från havets faror. Om du gör honom missnöjd riskerar du dina sjömäns liv."
"##new_festival##":"Anordna ny festival"
"##new_governor##":""
"##new_map##":"Fil"
"##new_trade_route_to##":"Ny handelsväg etablerad."
"##newcomer_this_month##":"nykomling anlände denna månad"
"##newcomers_this_month##":"nykomlingar anlände denna månad"
"##no_academy_access##":"Detta hus har inte tillgång till en högskola"
"##no_citizens_desire_live_here##":"Inga medborgare vill bo här"
"##no_culture_building_in_city##":"Du har ingen kultur i din stad, ergo (latin för därför) har du ingen kulturställning."
"##no_dock_for_sea_trade_routes##":"GLÖM INTE! Denna nya handelsrutt över havet kräver byggnation av en handelshamn innan några fartyg kan anlända."
"##no_fire_risk##":"Ingen brandrisk"
"##no_fishplace_in_city##":"Vår fiskebåt hoppas snart kunna hitta en fiskeplats. Det blir svårt att försörja sig om vi inte hittar fisk..."
"##no_food_stored_last_month##":"Inga livsmedel lagrades förra månaden"
"##no_goods_for_request##":"Du har inte tillräckligt med varor i dina handelsmagasin"
"##no_people_in_city##":"Inga människor i staden!"
"##no_priority##":"Ingen prioritet"
"##no_space_for_evolve##":"Denna boning skulle kunna få ännu högre status om den hade mer utrymme att expandera."
"##no_target_population##":"( Ingen målbefolkning )"
"##no_tax_in_this_year##":"Hittills i år har ingen skatt betalats från detta hus"
"##no_visited_by_taxman##":"Ej fått besök av skatteindrivare. Betalar ej skatt"
"##no_warning_for_us##":"Vi har inga rapporter om hot"
"##nomoney_for_gift_text##":"Du har inte tillräcklig med personliga besparingar för att kunna betala en gåva till kejsaren. Försök att betala dig själv högre lön!"
"##none_crime_risk##":"Ingen brottslighet i sikte här inte."
"##none_damage_risk##":"Ingen risk för kollaps"
"##northBtnTooltip##":""
"##not_available##":"Ej tillgänglig... ännu!"
"##not_need_education##":"Inga medborgare kräver ännu utbildningsmöjligheter. Men när staden börjar växa kommer människor att förvänta sig skolor och högskolor, och senare även bibliotek."
"##numidian_warrior##":"En numidisk soldat"
"##occupants##":"invånare"
"##oil_workshop_bad_work##":"Med så få anställda produceras nästan ingen olja alls. Det kommer mycket små leveranser av olja under det kommande året."
"##oil_workshop_full_work##":"Denna olivpress är fullt bemannad och producerar rikliga mängder olja av hög kvalitet."
"##oil_workshop_info##":"Här pressas olja från oliver, som plebejerna behöver för matlagning och för belysningen i sin Insulae. Överskottsoljan kan bli lönsam handel."
"##oil_workshop_need_resource##":"Denna olivpress kommer inte att producera olja utan leverans av oliver, från ett magasin eller från en lantgård."
"##oil_workshop_need_some_workers##":"Denna olivpress behöver fler arbetare för att nå sin fulla potential för oljeproduktion."
"##oil_workshop_no_workers##":"Denna olivpress har inga anställda och kommer inte att producera olja."
"##oil_workshop_no_workers##":"Detta krukmakeri har inga anställda. Produktionen har upphört."
"##oil_workshop_patrly_workers##":"Denna olivpress är underbemannad och producerar oljan mycket långsammare än vad den borde."
"##oil_workshop_slow_work##":"Mycket få människor arbetar vid denna olivpress. Som resultat är oljeproduktionen långsam."
"##oil_workshop##":"Oljepresseri"
"##oil##":"Olja"
"##ok##":"OK"
"##olive_factory_stock##":"Lagrade oliver,"
"##olive_farm_bad_work##":"De flesta träden har inga oliver eftersom nästan ingen arbetar här."
"##olive_farm_full_work##":"Denna lund har alla anställda den behöver. Trädgrenarna dignar med tunga lass av oliver."
"##olive_farm_info##":"Oliver är värdefulla för sin olja. Olivpresserierna ger olja för matlagning, belysning, smörjning och konservering."
"##olive_farm_need_some_workers##":"Denna lund utnyttjar inte maximal kapacitet. Olivproduktionen kan bli bättre med fler arbetare."
"##olive_farm_no_workers##":"Denna lantgård har inga anställda. Inget har planterats."
"##olive_farm_patrly_workers##":"Denna lund är underbemannad. Det tar längre tid att plocka oliverna än vad det borde."
"##olive_farm_slow_work##":"Det finns mycket få människor som arbetar här. Som resultat är olivproduktionen långsam."
"##olive_farm##":"Olivodling"
"##olive##":"Oliver"
"##open_trade_route##":"Öppna handelsväg"
"##options##":"Inställning"
"##oracle_info##":"Orakel ökar efterfrågan på husen i stadsdelen och gör de boende gladare. Denna byggnad tillfredsställer samtliga gudar."
"##oracle_need_2_cart_marble##":"Du behöver 2 ton marmor för att bygga ett orakel"
"##oracle##":"Orakel"
"##oracles_in_city##":"Orakel i staden"
"##oracles##":"Orakel"
"##other##":"Diverse"
"##our_foods_level_are_low##":"Våra livsmedelsförråd är små"
"##out_of_credit##":"Kredit saknas!"
"##overall_city_become_a_sleepy_province##":"Detta är på det hela taget en provins med få verkliga hot - precis så som invånarna vill ha det!"
"##overlays##":"Översikt"
"##ovrm_aborigen##":""
"##ovrm_academy##":""
"##ovrm_amphitheater##":"Amfiteatrar"
"##ovrm_barber##":""
"##ovrm_baths##":""
"##ovrm_clinic##":""
"##ovrm_colloseum##":""
"##ovrm_commerce##":""
"##ovrm_crime##":""
"##ovrm_damage##":""
"##ovrm_desirability##":""
"##ovrm_education##":"Allt"
"##ovrm_educations##":"Utbildning"
"##ovrm_entertainments##":""
"##ovrm_entrertainment##":"Allt"
"##ovrm_fire##":""
"##ovrm_food##":""
"##ovrm_health##":""
"##ovrm_hippodrome##":""
"##ovrm_hospital##":""
"##ovrm_library##":"Bibliotek"
"##ovrm_market##":"Marknadstillgång"
"##ovrm_religion##":""
"##ovrm_risks##":""
"##ovrm_school##":""
"##ovrm_simple##":""
"##ovrm_tax##":""
"##ovrm_text##":"Översikt"
"##ovrm_theater##":""
"##ovrm_tooltip##":""
"##ovrm_troubles##":""
"##ovrm_water##":""
"##partician_good_life##":"Var hälsad. Staden sköts riktigt bra."
"##partician_need_workers##":"Servicen blir lidande. Staden behöver fler arbetare."
"##patients#":"patienter"
"##patrician_average_life##":"Här i min bekväma villa anser jag livet i staden vara mycket bra."
"##patrician_gods_angry##":"Medborgare! Situationen är hotfull. Gudarna är vreda."
"##patrician_high_workless##":"Detta är skandalöst. Jag har aldrig sett så många arbetslösa plebejer."
"##patrician_low_entertainment##":"Medborgare! Är icke detta den tråkigaste staden i riket?"
"##patrician_so_hungry##":"Hell! Vad tjänar rikedom till om det inte finns mat att köpa?"
"##pay_to_open_trade_route?##":"Betala för att öppna denna väg?"
"##peace_rating_text##":"Fredsställningen blir bättre för varje år utan upplopp eller invasioner som skadar egendom i städerna."
"##peaceful_crime_risk##":"Detta är en fridfull stadsdel."
"##people_leave_city_insane_tax##":"Människor lämnar staden på grund av dina höga skatter"
"##people_leave_city_low_wage##":"Människor beger sig av på jakt efter högre löner"
"##people_leave_city_some##":"Människor lämnar staden"
"##people##":"denarer"
"##percents##":"Ränta på"
"##person##":"denarer"
"##plaza_caption##":"Torg"
"##plaza##":"Torg"
"##plname_continue##":"Fortsätt"
"##plname_start_new_game##":"Ny karriär"
"##pn_salary##":"Personlig inkomst"
"##poor_city_mood_lack_migration##":"Stämningen i staden förhindrar immigration"
"##poor_housing_discourages_migration##":"Dåliga bostäder motverkar invandring trots välståndet i staden"
"##pop##":"Inv"
"##population_registered_as_taxpayers##":"av befolkningen är skatteskrivna"
"##population_tooltip##":"Befolkningsmängd"
"##population##":"Befolkning"
"##pottery_bad_work##":"Mycket få människor arbetar här. Som resultat går krukproduktionen långsamt."
"##pottery_workshop_bad_work##":"Med så få anställda vid krukmakeriet står produktionen nästan stilla. Det kommer inte att produceras mycket krukor under det kommande året."
"##pottery_workshop_full_work##":"Detta krukmakeri har alla anställda det behöver. Det arbetar fullt ut med att producera krukor."
"##pottery_workshop_info##":"Här formar krukmakare lera till kärl som medborgarna använder till förvaring. Handla med krukor, eller låt dina marknader distribuera dem så att människorna kan bygga bättre hus."
"##pottery_workshop_need_resource##":"Detta krukmakeri behöver leveranser av lera, från ett magasin eller från ett lertag, för att kunna producera krukor."
"##pottery_workshop_need_som_workers##":"Detta krukmakeri är underbemannat och produktionen tar längre tid än normalt."
"##pottery_workshop_patrly_workers##":"Detta krukmakeri utnyttjar inte maximal kapacitet. Som resultat kommer krukproduktionen att gå långsammare."
"##pottery_workshop##":"Krukmakeri"
"##pottery##":"Krukor"
"##praetor_salary##":"Pretorslön på"
"##prefect_fight_fire##":"Hettan från elden är otroligt stark."
"##prefect_gods_angry##":"Jag är rädd för att gudarna kommer att förbanna staden."
"##prefect_good_life##":"Detta är en underbar plats att bo på."
"##prefect_high_workless##":"Jag har aldrig sett så många arbetslösa!"
"##prefect_high_workless##":""
"##prefect_low_entertainment##":"Brottslingarna jag tar får bättre underhållning än den här staden!"
"##prefect_need_workers##":"Denna stad är i desperat behov av arbetare!"
"##prefect_so_hungry##":"Det finns inte nog med mat i staden. Det ökar brottsligheten."
"##prefecture_bad_work##":"Vi arbetar endast med kontorspersonal. Det går ofta en hel månad utan att vi sänder en prefekt ut på gatorna."
"##prefecture_full_work##":"För närvarande är vår tjänstgöringslista full. Våra prefekter är alltid ute och patrullerar gatorna."
"##prefecture_info##":"Prefekturerna sänder prefekter till staden för att hålla fred, och för att bekämpa bränder. Ordning kan endast upprätthållas om prefekterna patrullerar staden."
"##prefecture_need_some_workers##":"Vi har lite ont om prefekter. Vi har luckor på en dag eller två i vår täckning."
"##prefecture_no_workers##":"Utan personal blir den här stationen inte mycket mer än en måltavla för vandaler."
"##prefecture_on_patrol##":"Vår prefekt är ute och patrullerar."
"##prefecture_patrly_workers##":"Vi är underbemannade, och har farliga luckor på upp till en vecka i vår tjänstgöringslista."
"##prefecture_ready_for_work##":"Vår prefekt förbereder sig för sin tjänst."
"##prefecture_slow_work##":"Vi har alldeles för få prefekter. Det händer att inga prefekter lämnar stationen på upp till två veckor åt gången."
"##prefecture##":"Prefektur"
"##prepare_to_festival##":"Förbereder den kommande festivalen"
"##press_escape_to_exit##":"Högerklicka för att avsluta"
"##priest_gods_angry##":"Vi är i fara! Staden visar ingen respekt för gudarna."
"##priest_good_life##":"Livet är mycket behagligt i denna stad."
"##priest_good_life##":"Denna stad är en hygglig plats att bo på."
"##priest_high_workless##":"Arbetslösheten är oroväckande hög."
"##priest_low_entertainment##":"Denna stad är så tråkig. Även en präst tycker om gladiatorspel då och då."
"##priest_need_workers##":"Detta ställe behöver många fler arbetare."
"##priest_so_hungry##":"Var hälsad. Denna stad behöver omedelbart mer livsmedel."
"##priority_button_tolltip##":"Klicka på ett nummer för att fastställa prioritetsnivå. Alla övriga uppgifter kommer att omjusteras"
"##priority_level##":"Prioritetsnivå"
"##proconsoul_salary##":"Prokonsulslön på"
"##procurator_salary##":"Prokuratorslön på"
"##profit##":"Nettoflöde in/ut"
"##prosperity_lack_that_you_pay_less_rome##":"Att betala lägre löner än Rom ger din stad rykte att vara mindre blomstrande."
"##province_has_peace_a_short_time##":"Denna provins har haft fred en kort tid, men dina invånare känner sig fortfarande inte helt säkra. Fler fredsår kommer att förbättra detta."
"##qty_stacked_in_city_warehouse##":"i handelsmagasin"
"##quaestor_salary##":"Kvestorslön på"
"##quarry_bad_work##":"Det finns nästan inga anställda vid det här brottet, och produktionen står nästan stilla."
"##quarry_full_work##":"Detta brott har alla anställda det behöver, det arbetar fullt ut med att producera marmor."
"##quarry_info##":"Bryt marmor ur intilliggande klippor och använd den till att bygga orakel och stora tempel. Marmor är vanligen en värdefull exportvara."
"##quarry_need_some_workers##":"Detta brott utnyttjar inte maximal kapacitet. Som resultat kommer marmorproduktionen att bli något mindre."
"##quarry_no_workers##":"Detta brott har inga anställda. Produktionen har upphört."
"##quarry_patrly_workers##":"Mycket få människor arbetar vid det här brottet. Som resultat är marmorproduktionen långsam."
"##quarry_slow_work##":"Mycket få människor arbetar vid detta lertag. Som resultat är lerproduktionen långsam."
"##quarry##":"Marmorbrott"
"##quit##":"Avsluta"
"##rating##":"Ställning"
"##rawm_production_complete_m##":"Produktionen är"
"##ready_to_game##":""
"##really_destroy_fort##":"Är du säker på att du vill ta detta fort ur aktiv tjänst?"
"##recruter_gods_angry7##":"Vi har problem! Gudarna är förargade på oss."
"##recruter_good_life##":"Var hälsad! Livet här är gott."
"##recruter_high_workless##":"Var hälsad! Har du sett hur hög arbetslösheten är?"
"##recruter_low_entertainment##":"Jag arbetar hårt och jag vill roa mig ofta. Men det går inte här. Det finns inget att göra!"
"##recruter_need_workers##":"Medborgare! Denna stad behöver fler arbetare."
"##recruter_normal_life##":"Var hälsad. Detta är en ganska bra stad."
"##recruter_so_hungry##":"Kan du avvara lite bröd? Jag har inte ätit på så länge."
"##reject##":"Avvisa varor"
"##religion_access_1_temple##":"Detta hus har endast tillgång till ett tempel för en enda gud"
"##religion_access_2_temple##":"Detta hus har tillgång till tempel för 2 olika gudar"
"##religion_access_3_temple##":"Detta hus har tillgång till tempel för 3 olika gudar"
"##religion_access_4_temple##":"Detta hus har tillgång till tempel för 4 olika gudar"
"##religion_access_5_temple##":"Detta hus har tillgång till tempel för alla gudarna"
"##religion_access_full##":"Detta hus har tillgång till ett orakel, och till tempel för alla gudar"
"##religion_advisor##":"Religiösa byggnader"
"##religion_in_your_city_is_flourishing##":"Religionen i din stad blomstrar. Invånarnas olika religionsbehov uppfylls, och prästerna rapporterar att gudarna är nöjda."
"##religion_no_access##":"Detta hus har inte tillgång till några tempel eller orakel"
"##religion##":"Religion"
"##religionadv_need_basic_religion##":"Fler och fler medborgare kräver minst en gudstjänstplats i sitt bostadsområde, för att förbättra gudarnas uppfattning om dem."
"##religionadv_need_second_religion##":"Medborgarna i vissa områden vill ha tillgång till en annan religion nära hemmet. Bristen på religioner hindrar stadens utveckling i vissa områden."
"##religionadv_need_third_religion##":"Vissa medborgare vill ha en tredje religion etablerad nära sitt område. De anser att detta skulle attrahera bättre patricierklasser."
"##replay_game##":"Börja om"
"##request_btn_tooltip##":"Klicka här för att sända iväg begäran"
"##request_failed##":"Din nyligen visade oförmåga eller ovilja att utföra en kejserlig begäran har skadat din ställning i Rom en aning."
"##requierd##":"Behov"
"##reservoir_info##":"Denna gigantiska cistern innehåller rent dricksvatten, som distribueras via rör av lera över en stor radie i staden. Akvedukter kan länka samman reservoarerna över stora avstånd."
"##reservoir_no_water##":"Denna reservoar fungerar inte eftersom den inte ligger intill vatten eller inte är ansluten till en annan reservoar via akvedukter."
"##reservoir##":""
"##restocking_fishing_boat##":"Vi förbereder för närvarande vår fiskebåt för att segla ut igen. Hur snabbt det går beror på hur många anställda vi har."
"##return_2_fort##":"Återvänd till fortet"
"##return_to_main_map##":"Återvänd till spelets huvudkarta"
"##rift_info##":"Sprickor i marken"
"##right_click_to_exit##":"Högerklicka för att avsluta"
"##rioter_say_1##":"Ståthållaren bryr sig uppenbarligen inte om mig, så jag tänker visa vad jag tycker om hans stad."
"##rioter_say_3##":"Om du vill veta hur städer ser ut när de brinner, se noga på nu!"
"##rladv_mood##":"Gudarna är"
"##road_caption##":"Väg"
"##road_from_rome##":"Detta är vägen till Rom. Immigranterna anländer från denna punkt. Därför är det viktigt att vägen hålls öppen. Även köpmän passerar genom din provins längs denna kejserliga huvudväg."
"##road_text##":"Vägarna är livsviktiga för stadens funktion. Invånarna går bara ut ur sina hus om det finns en väg."
"##road_to_distant_region##":"Detta är den väg som leder till rikets utposter. Det är en kejserlig huvudväg, som måste hållas öppen längs hela sin sträckning."
"##roadBtnTooltip##":""
"##rock_caption##":"Klippor"
"##rock_text##":"Klipporna kan inte forceras eller röjas undan. Marmor- och malmbrott fungerar bara om de uppförs nära klippor."
"##roman_city##":"En romersk stad"
"##rome_prices##":"Priser fastställs av Rom"
"##romeGuard_average_life##":"Allt verkar lugnt här."
"##romeGuard_gods_angry##":"Gudarna är förargade på denna plats."
"##romeGuard_good_live##":"Jag må vara en simpel soldat, men även jag kan se vilken storslagen stad detta är."
"##romeGuard_high_workless##":"I dessa tider av arbetslöshet tackar jag gudarna att jag har jobb."
"##romeGuard_low_entertainment##":"Om det fanns bättre underhållning i staden skulle vakttjänsten inte kännas så betungande."
"##romeGuard_need_workers##":"Den här staden behöver många fler arbetare."
"##romeGuard_so_hungry##":"Hur ska en soldat kunna slåss utan mat?"
"##rotateLeftBtnTooltip##":""
"##rotateRightBtnTooltip##":""
"##samnite_soldier##":"En samnitisk soldat"
"##save_city##":"Spara spel"
"##save_game_here##":"Spara det aktuella spelet till denna fil"
"##save_map##":"Öppna karta"
"##scholar_average_life##":"Den här staden verkar bra."
"##scholar_gods_angry##":"Hjälp! Gudarna är vreda. De kommer att straffa oss."
"##scholar_good_life##":"Den här staden är fantastisk."
"##scholar_high_workless##":"Det är jättemånga som söker arbete här."
"##scholar_low_entertainment##":"Staden är så tråkig. Jag vill se fler föreställningar."
"##scholar_need_workers##":"Det finns så få arbetare att någon till och med erbjöd mig jobb."
"##scholar_so_hungry##":"Jag svälter ihjäl!"
"##scholar##":"Skolbarn"
"##scholars##":"i skolålder"
"##school_access_perfectly##":"Områden som kräver utbildningsmöjligheter har tillgång till dem, men fler skolor skulle minska storleken på klasserna."
"##school_full_access##":"Detta hus har tillgång till skola"
"##school_full_work##":"Denna skola används, och barnen i stadsdelen är läskunniga och vältaliga."
"##school_info##":"Barn måste gå i stadsdelsskolorna för att lära sig grunderna i läsning, skrivning och retorik om de skall kunna växa upp till produktiva vuxna."
"##school_no_access##":"Detta hus har inte tillgång till någon skola"
"##school_no_workers##":"Denna skola används inte, och är värdelös för lokalsamhället."
"##school##":"Skola"
"##schools##":"Skolor"
"##screen_settings##":"Bild"
"##scribe_messages_title##":"Meddelanden från dina skrivare"
"##scribemessages_unread##":"Oläst meddelande. Vänsterklicka på detta meddelande för att läsa det.  Högerklicka på detta meddelande för att radera det"
"##scrw_subject##":"Ämne"
"##sdlr_bold##":"Modig"
"##seamerchant_noany_trade##":"Om jag fick bestämma skulle jag inte segla den här vägen. Den här staden varken köper eller säljer något."
"##select_city_layer##":"Välj en översiktsrapport för staden"
"##select_location##":""
"##seleucid_soldier##":"En selucidisk soldat"
"##sell_price##":"Säljarna får"
"##senate_1_info##":"Senatsbyggnaden är en av de attraktivaste byggnaderna i staden. Den ger anställning åt skatteindrivarna och inkomsterna från deras verksamhet förvaras här."
"##senate_1##":"Senat"
"##senate_save##":"i stadskassan"
"##senate##":"Senat"
"##senateBtnTooltip##":""
"##senatepp_clt_rating##":"Kultur"
"##senatepp_favour_rating##":"Popularitet"
"##senatepp_peace_rating##":"Fred"
"##senatepp_prsp_rating##":"Välstånd"
"##senatepp_unemployment##":"Arbetslöshet"
"##send_generous_gift##":"Sänd en generös gåva"
"##send_lavish_gift##":"Sänd en frikostig gåva"
"##send_legion_to_emperor##":"Be din militära rådgivare att avdela några stridsklara legioner i imperiets tjänst"
"##send_modest_gift##":"Sänd en blygsam gåva"
"##send_money_to_city##":"Ge pengar till staden"
"##send_money##":"Donera dessa pengar till staden från dina personliga besparingar"
"##send_to_city##":"Ge till staden"
"##sentiment_people_angry_you##":"Människorna är arga på dig"
"##sentiment_people_annoyed_you##":"Människorna är förargade på dig"
"##sentiment_people_extr_pleased_you##":"Människorna är extremt nöjda med dig"
"##sentiment_people_idolize_you##":"Människorna avgudar dig, som en gud"
"##sentiment_people_indiffirent_you##":"Människorna är likgiltiga inför dig"
"##sentiment_people_love_you##":"Människorna älskar dig"
"##sentiment_people_pleased_you##":"Människorna är nöjda med dig"
"##sentiment_people_upset_you##":"Människorna är upprörda över dig"
"##sentiment_people_veryangry_you##":"Människorna är mycket arga på dig"
"##sentiment_people_verypleased_you##":"Människorna är mycket nöjda med dig"
"##sentiment_people_veryupset_you##":"Människorna är mycket upprörda över dig"
"##set_amount_to_donate##":"Fastställ summa att donera"
"##set_mayor_salary##":"Klicka här för att fastställa din personliga lön"
"##several_crimes_but_area_secure##":"Flera brott har rapporterats här nyligen, men på det hela taget har prefekterna situationen under kontroll"
"##shipyard_info##":"Med några vagnslaster timmer och tillräckligt med arbetare bygger fartygsvarvet fiskebåtar till stadens fiskehamnar."
"##shipyard_notneed_ours_boat##":"Det finns för närvarande inga fiskehamnar som behöver våra båtar."
"##shipyard##":"Fartygsvarv"
"##show_bigpanel##":"Visa hela sidopanelen"
"##show_prices##":"Visa priser"
"##show_spots_of_city_troubles_tip##":"Växla mellan aktuella problemområden i staden"
"##show##":"Evenemang"
"##showing_agamemnon_aeschylus##":"Uppför: 'Annales', av Tacitus"
"##showing_antigone_sophocles##":"Uppför: Homeros grekiska tragedier"
"##showing_lisistrata_aristopanes##":"Uppför: 'Vergilius dikter'"
"##showing_odyssey_homer##":"Uppför: 'Platons filosofi'"
"##showing_thecrito_plato##":"Uppför: 'Oidipus', av Sofokles"
"##simple_formation_text##":"En enkel formation, som ger fördelar åt försvarstrupper."
"##sldh_health_sparse##":"Gles"
"##sldh_health_strong##":"Stark"
"##sldh_health_strongest##":"Extremt stark"
"##sldr_badly_shaken##":"Mycket uppskakad"
"##sldr_daring##":"Djärv"
"##sldr_encouraged##":"Uppmuntrad"
"##sldr_extremely_scared##":"Extremt rädd"
"##sldr_shaken##":"Uppskakad"
"##sldr_terrified##":"Livrädd"
"##sldr_totally_distraught##":"Vettskrämd"
"##sldr_very_bold##":"Mycket modig"
"##sldr_very_frightened##":"Mycket rädd"
"##small_ceres_temple##":"Cerestempel"
"##small_colloseum_show##":"Det krävs fler spektakel i dina colosseum! Genom att förse dem med gladiatorer eller lejon förbättras underhållningen i delar av staden."
"##small_domus##":"Liten Insulae"
"##small_festival##":"Liten festival"
"##small_food_on_next_month##":"- mycket lite mat kommande månad"
"##small_hovel##":"Litet skjul"
"##small_hut##":"Litet hus"
"##small_mars_temple##":"Marstempel"
"##small_mercury_temple_info##":"Handelsmännen dyrkar Merkurius för att skydda sina varor. Om Merkurius vrede väcks sätts allas vinst på spel."
"##small_mercury_temple##":"Merkuriustempel"
"##small_neptune_temple##":"Neptunustempel"
"##small_palace##":"Litet palats"
"##small_shack##":"Liten koja"
"##small_temples##":"Små tempel"
"##small_tent##":"Litet tält"
"##small_venus_temple##":"Venustempel"
"##small_villa##":"Liten villa"
"##small##":"Litet"
"##smallcurse_of_mars_text##":"Mars, soldaternas beskyddare och segerförlänare, är missnöjd. Dina soldater fruktar att de kommer att förlora ett stort slag om han inte blidkas."
"##smallcurse_of_mercury_description##":"Merkurius, gudarnas budbärare och handelsmännens beskyddare, är missnöjd. Dina handelsmän fruktar att hans beskydd viker."
"##smcurse_of_venus_description##":"Venus, förmedlare av kärlek och harmoni, är upprörd. Detta bådar inget gott för prefekterna i din stad!"
"##smcurse2_of_venus_description##":"När Venus är missnöjd sänker hon medborgarnas sinnesstämning. En del säger att hon för med sig sjukdomar."
"##soldier##":"Soldat"
"##soldiers_health##":"Soldaternas hälsa"
"##soldiers_in_legion##":"Soldater i legion"
"##soldiers##":"Soldater"
"##some_amphitheaters_no_actors##":"Vissa av dina amfiteatrar saknar skådespelare och gladiatorer. Fler underhållare skulle ge bättre villkor i de stadsdelar som klagar över dålig underhållning."
"##some_crime_risk##":"Området löper viss risk att drabbas av brottslighet."
"##some_defects_damage_risk##":"Mycket liten risk för kollaps"
"##some_fire_risk##":"Viss brandrisk"
"##some_food_on_next_month##":"- vissa livsmedel kommande månad"
"##some_houses_inadequate_entertainment##":"Vissa medborgare klagar över bristande tillgång till underhållning i sina områden. Du kanske behöver erbjuda ett mer varierat utbud, eller kanske bygga fler skådespelarkolonier till dina teatrar."
"##some_houses_need_amph_for_grow##":"Vissa medborgare klagar över bristande tillgång till fritidsanläggningar. Vissa områden i staden kräver mer varierade underhållningsmöjligheter."
"##some_houses_need_better_library_access##":"Vissa områden i staden vill ha bättre tillgång till bibliotek. Välbärgade medborgare tycker om att läsa men vill inte gå långt för att nå biblioteket."
"##some_houses_need_library_or_colege_access##":"Vissa områden i staden kräver nu skolor och högskolor. Bristen på utbildningsmöjligheter förhindrar byggandet av bättre bostäder i dessa områden."
"##some_low_fire_risk##":"Denna byggnad utgör en försumbar brandrisk"
"##sound_settings##":"Ljud"
"##spear##":"Spjut"
"##special_orders##":""
"##speed_settings##":"Hastighet"
"##spirit_of_mars_text##":""
"##spirit_of_mars_title##":""
"##stacking_resource##":"Hamstrar vara"
"##stacking##":"Hamstrar"
"##start_condition##":"Startvillkor"
"##start_this_map##":""
"##statue_big_info##":"Monument över framstående medborgare och historiska händelser ger ett område bättre status. Folket är stolta över att ha statyer i grannskapet... och ju större desto bättre."
"##statue_big##":"Stor staty"
"##statue_desc##":""
"##statue_middle##":"Medelstor staty"
"##status_small##":"Liten staty"
"##stop_granary_devastation##":"Sluta tömma sädesmagasin"
"##stop_warehouse_devastation##":"SLUTA tömma magasin"
"##students##":"i högskoleålder."
"##syracusae_somewhat_dangerous_province##":"Syracusae: en något farlig provins"
"##tamer_normal_life##":"Om du rör mitt lejon, får du smaka på min piska."
"##tarentum_slightly_dangerous_province##":"Tarentum: en inte helt ofarlig provins"
"##tarentum_win_text##":"Etruskerna kommer inte att hota Tarentum igen. Bra gjort! Det är sällsynt med en ståthållare som finner rätt balans mellan stadsbyggnation och strid. Låt se om du kan göra om din bravad eller om det bara handlade om tur."
"##target_population_is##":"( Målbefolkningen är"
"##tarraco_peaceful_province##":"Tarraco: en fredlig provins"
"##tarraco_win_text##":"Tarracos livsmedelsexport hjälpte imperiet att överleva en svår period. Medborgarna är skyldiga dig för sina liv och ståthållarna sina arbeten. Skördarna blir nu normala igen och jag vill använda dina talanger inom ett nytt område."
"##tarsus_largerly_peacefull_province##":"Tarsus: en mestadels fredlig provins"
"##tarsus_win_text##":"Du är på god väg att bli min mest uppskattade undersåte. Din mästerliga förståelse av handeln gjorde Tarsus till precis den stad jag hoppats på. De östliga provinserna är mer lojala i dag, tack vare dig."
"##tax_rate##":"Skattesatsen"
"##taxCollector_average_life##":"Staden tycks fungera väl."
"##taxCollector_gods_angry##":"Om vi inte bygger fler tempel snart, kommer gudarna att förbanna denna stad."
"##taxCollector_good_life##":"Var hälsad! Detta är en mycket trevlig stad att bo i."
"##taxCollector_high_tax##":"Har du sett skatterna här? Medborgare, det är inte rätt."
"##taxCollector_high_workless##":"Jag ogillar det här stället. Arbetslösheten är för hög."
"##taxCollector_low_entertainment##":"Jag skulle inte ha nåt emot att pressa folk på denarer hela dagarna om det bara fanns mer att göra på kvällarna!"
"##taxCollector_need_workers##":"Den här staden behöver fler arbetare och det genast."
"##taxCollector_so_hungry##":"Om vi inte får mer livsmedel finns det snart ingen som kan betala skatt!"
"##taxCollector_very_little_tax##":"Dessa hus betalar så lite skatt att det är slöseri med tiden."
"##taxes##":"Inkasserade skatter"
"##taxСollector_low_tax_collected##":"Att driva in skatt från dessa hårt arbetande människor får mig nästan att gråta - men bara nästan!"
"##taxСollector_much_tax##":"Jag älskar att driva in skatt från rika hus som dessa."
"##teacher_average_life##":"Jag ger staden åtta av tio poäng."
"##teacher_gods_angry##":"Vi får känna gudarnas vrede om vi inte bygger fler tempel snart."
"##teacher_good_life##":"Staden får full pott. Det är en underbar plats."
"##teacher_high_workless##":"Bara jag inte förlorar jobbet. Arbetslösheten är så hög att jag inte skulle få ett nytt."
"##teacher_low_entertainment##":"Staden är så tråkig! Den behöver mer underhållning."
"##teacher_need_workers##":"Otroligt att det finns så många arbetstillfällen här."
"##teacher_so_hungry##":"Det saknas livsmedel här. Det gör medborgarna olyckliga."
"##templeBtnTooltip##":""
"##temples##":"Tempel"
"##testers##":""
"##thanks_to##":""
"##theater_full_access##":"Detta hus har tillgång till teater"
"##theater_full_work##":"Denna teater sätter för närvarande upp pjäser med lokala aktörer, som vanligen drar stor publik."
"##theater_need_actors##":"Teatrarna och amfiteatrarna söker alltid efter nya talanger."
"##theater_no_access##":"Detta hus har inte tillgång till en teater"
"##theater_no_have_any_shows##":"Denna teater har sällan några uppsättningar. Den behöver riktiga skådespelare för att kunna erbjuda underhållning."
"##theater_no_workers##":"Vinden är det enda som rör sig i denna teater. Utan arbetare erbjuder den inga pjäser till lokalbefolkningen."
"##theater##":"Teater"
"##theaters##":"Teatrar"
"##these_rift_info##":"Dessa klyftor har orsakats av jordbävningar. De kan inte passeras eller fyllas."
"##this_fire_can_spread##":"Dessa eldsvådor sprider sig om du inte snabbt hejdar dem."
"##this_is_ruins##":"Detta är spillrorna från byggnaden som nämns ovan. Förfallna platser gör inte att området ser vackrare ut."
"##this_lawab_province_become_very_peacefull##":"Detta är en laglydig provins som med tiden kan bli mycket fredlig."
"##this_time_you_city_not_need_religion##":"Dina medborgare är ännu så länge upptagna med andra aspekter på stadslivet. I takt med att staden växer kommer de att vilja ha tillgång till ett stort Tempelutbud."
"##this_year##":"Så här långt detta året"
"##timber_factory_stock##":"Lagrat virke,"
"##timber_mill_need_trees##":"Bygg brädgård intill träden"
"##timber##":"Timmer"
"##time_since_last_gift##":"Tid sedan senaste gåva"
"##tingis_dangerous_province##":"Tingis: en farlig provins"
"##tingis_win_text##":"Är du ståthållare eller general? Din utmärkta insats vid Tingis befriar mina legioner från tjänstgöring i väst och låter mig ägna tiden åt andra strävanden. Du börjar bli en nyckelperson i min planering."
"##to_empire_road##":"Till Imperiet"
"##to_rome_road##":"Till Rom"
"##to_trade_advisor##":"Till handelsrådgivaren"
"##tooltip_full##":"Mushjälp FULL"
"##tooltip_some##":"Mushjälp HALV"
"##tower_have_workers_no_soldiers##":"Vi har underhållspersonal, men vi behöver trupper från en förläggning för att försvara staden."
"##tower_may_build_on_thick_walls##":"Du kan endast bygga torn på tjocka murar"
"##tower_need_wall_for_patrol##":"Måste finnas intill en mur för att sända ut en patrull"
"##tower_no_workers##":"Utan bemanning har vi ingen personal till våra kastmaskiner eller vakter som kan patrullera murarna."
"##tower##":"Torn"
"##trade_advisor_blocked_clay_production##":"Din handelsrådgivare har stoppat alla lertag."
"##trade_advisor_blocked_fruit_production##":"Din handelsrådgivare har stoppat all fruktodling."
"##trade_advisor_blocked_furniture_production##":"Din handelsrådgivare har stoppat all möbeltillverkning."
"##trade_advisor_blocked_grape_production##":"Din handelsrådgivare har stoppat all druvodling."
"##trade_advisor_blocked_iron_production##":"Din handelsrådgivare har stoppat all malmbrytning."
"##trade_advisor_blocked_marble_production##":"Din handelsrådgivare har stoppat all marmorbrytning."
"##trade_advisor_blocked_meat_production##":"Din handelsrådgivare har stoppat all köttproduktion."
"##trade_advisor_blocked_oil_production##":"Din handelsrådgivare har stoppat all oljeproduktion."
"##trade_advisor_blocked_olive_production##":"Din handelsrådgivare har stoppat all olivodling."
"##trade_advisor_blocked_pottery_production##":"Din handelsrådgivare har stoppat all kruktillverkning."
"##trade_advisor_blocked_timber_production##":"Din handelsrådgivare har stoppat all avverkning."
"##trade_advisor_blocked_vegetable_production##":"Din handelsrådgivare har stoppat all grönsaksodling."
"##trade_advisor_blocked_weapon_production##":"Din handelsrådgivare har stoppat all vapenproduktion."
"##trade_advisor_blocked_wheat_production##":"Din handelsrådgivare har stoppat all veteodling."
"##trade_advisor_blocked_wine_production##":"Din handelsrådgivare har stoppat all vinproduktion."
"##trade_advisor##":"Handelsrådgivare"
"##trade_btn_notrade_text##":"Gör ej affärer"
"##trade_caravan_from##":"Köpmannakaravan från"
"##trade##":"Handel"
"##tradeadv_industrystate_tip##":"Starta eller avsluta produktion för denna aktivitet överallt i staden"
"##trees_and_forest_caption##":"Träd och skogsland"
"##trees_and_forest_text##":"Träden kan inte forceras, men de kan röjas undan. De är livsviktiga för skogsindustrin, brädgårdar måste ligga nära träden för att producera timmer."
"##triumphal_arch_info##":"Detta magnifika byggnadsverk är tillägnat Roms historiska segrar över sina fiender. Inget kan ge högre status."
"##triumphal_arch##":"Triumfbåge"
"##trouble_colloseum_full_work##":"Detta colosseum har både gladiatorkamp och lejonkamper, till lokalsamhällets stora nöje."
"##trouble_colloseum_have_only_gladiatros##":"Detta colosseum har gladiatorkamp för lokalbefolkningen. Lejon skulle ge mer variation till dödskamperna."
"##trouble_colloseum_have_only_lions##":"Detta colosseum har djurkamp, med lejon från lokala handelsmän. Den skulle också kunna anlita gladiatorer för kamp man mot man."
"##trouble_colloseum_no_shows##":"Detta colosseum ger inga föreställningar. Det behöver gladiatorer och lejon för att attrahera publik."
"##trouble_farm_was_blighted_by_locust##":"Jordbrukets marker har skadats av gräshoppssvärmarna, återhämtningen kommer att ta tid."
"##trouble_have_damage##":"Denna byggnad löper en liten risk att kollapsa"
"##trouble_hippodrome_full_work##":"Denna hippodrom har ofta spännande kapplöpningar, som ger mycket nöje åt lokalbefolkningen."
"##trouble_hippodrome_no_charioters##":"Denna hippodrom kör inga kapplöpningar. Den behöver körsvenner."
"##trouble_low_fire_risk##":"Denna byggnad har ingen brandrisk"
"##trouble_most_damage##":"Denna byggnad har många strukturella brister och sprickor"
"##trouble_most_fire##":"Denna byggnad är en brandfara"
"##trouble_need_olive##":"Denna byggnad kräver oliver"
"##trouble_need_road_access##":"Denna byggnad kräver åtkomst till väg"
"##trouble_need_timber##":"Denna byggnad kräver timmer"
"##trouble_no_damage##":"Denna byggnad är i perfekt strukturellt skick"
"##trouble_some_damage##":"Denna byggnad löper försumbar risk att kollapsa"
"##trouble_some_fire##":"Denna byggnad har brandrisk"
"##trouble_too_far_from_water##":"Denna byggnad är inte intill vatten!"
"##try_reduce_your_high_salary##":"Rom tycker att din lön är för hög för din nuvarande ställning. Du borde sänka den lite."
"##try_reduce_your_salary##":"Rom tycker att din lön är för hög för din nuvarande ställning. Det skulle vara bra om du sänkte den."
"##tutorial_prefecture_info##":""
"##tutorial_win_text##":"Gratulerar! Du har förstått grunderna på ett nöjsamt sätt. För att på bästa sätt fortsätta din utbildning, har jag ännu ett lindrigt uppdrag åt dig. Mot Brundisium!"
"##tutorial2_win_text##":"Du lär dig snabbt! Nu har du tillräckligt med kunskap för att klara ett riktigt uppdrag. Från och med nu kan du välja vilken riktning din karriär ska ta. Välj en fredligare provins om du vill koncentrera dig på att styra eller en farligare provins om du vill tampas med Roms fiender."
"##unable_fullfill_request##":"Kan inte fullgöra begäran"
"##unit##":"År"
"##units_in_stock##":"Lagrar"
"##units##":"År"
"##use_and_trade_resource##":"Använder och byteshandlar med denna vara"
"##valencia_peacefully_province##":"Valentia: en relativt fredlig provins"
"##valencia_win_text##":"Hispaniens nya huvudstad är precis vad vi behöver för att knyta den avlägsna provinsen tätare till Rom. Genom att krossa etruskerna så totalt försvinner det sista hotet i väst."
"##valentia_preview_mission##":"Ståthållaren ställs inför olika hot och faror, och Iberierna utgör inte det minsta av dessa! De har inte för avsikt att ge upp Hispanien."
"##vegetable_farm_bad_work##":"Det finns knappt några anställda för att underhålla jordbruket, de få grönsakerna kommer att bli offer för insekter."
"##vegetable_farm_full_work##":"Denna lantgård har alla anställda det behöver. Grönsaker växer här i överflöd."
"##vegetable_farm_info##":"Grönsaker är en viktig del av den balanserad diet som ditt folk behöver för hälsa och glädje. I sädesmagasinen lagras grönsaker för lokal konsumtion, och i handelsmagasinen förvaras överskottet för export."
"##vegetable_farm_need_some_workers##":"Denna lantgård är underbemannad. Vissa av dess grönsaker kommer att ruttna på åkern."
"##vegetable_farm_no_workers##":"Denna lantgård har inga anställda. Inget har planterats."
"##vegetable_farm_no_workers##":"Denna lund har inga anställda. Produktionen har upphört."
"##vegetable_farm_patrly_workers##":"Denna lantgård utnyttjar inte maximal kapacitet. Därför kommer grönsaksproduktionen att gå något långsammare."
"##vegetable_farm_slow_work##":"Mycket få jordbrukare arbetar här. De få grönsaker som odlas är små och osunda."
"##vegetable_farm##":"Grönsaksodling"
"##vegetable##":"Grönsaker"
"##venus_desc##":"Kärlek"
"##venus##":"Venus"
"##very_high_damage_risk##":"Denna byggnad är ostadig, och kommer sannolikt att falla samman snart"
"##very_high_fire_risk##":"Mycket stor brandrisk"
"##very_low_crime_risk##":"Detta är en mycket laglydig stadsdel, ingen brottslighet alls"
"##very_low_damage_risk##":"Denna byggnad har vissa strukturella brister"
"##very_low_fire_risk##":"Mycket liten brandrisk"
"##vinard_bad_work##":"Det finns mycket få anställda på denna odling. Som resultat kommer mycket få druvor att klara sig till skörden."
"##vinard_full_work##":"Denna odling har alla anställda den behöver. Vinrankorna är tunga med stora, saftiga druvor."
"##vinard_info##":"Druvorna från dessa vinrankor har odlats särskild för vinframställning. Vingårdarna gör fint vin för dina egna patricier, samt för export."
"##vinard_need_some_workers##":"Denna odling är underbemannad. Det tar längre tid att producera druvor än vad det borde."
"##vinard_no_workers##":"Denna odling har inga anställda. Produktionen har upphört."
"##vinard_patrly_workers##":"Denna odling utnyttjar inte maximal kapacitet. Som resultat kommer druvproduktionen att bli mindre."
"##vinard_slow_work##":"Mycket få människor arbetar på denna odling. Som resultat är druvproduktionen långsam."
"##vinard##":"Druvodling"
"##vinard##":"Vindruvsodling"
"##visit_chief_advisor##":"Besök din huvudrådgivare"
"##visit_education_advisor##":"Besök din utbildningsrådgivare"
"##visit_entertainment_advisor##":"Besök din underhållningsrådgivare"
"##visit_financial_advisor##":"Besök din finansrådgivare"
"##visit_health_advisor##":"Besök din hälsorådgivare"
"##visit_imperial_advisor##":"Besök din imperierådgivare"
"##visit_labor_advisor##":"Besök din arbetsrådgivare"
"##visit_military_advisor##":"Besök din militärrådgivare"
"##visit_population_advisor##":"Besök din befolkningsrådgivare"
"##visit_rating_advisor##":"Besök din ställningsrådgivare"
"##visit_religion_advisor##":"Besök din religionsrådgivare"
"##visit_trade_advisor##":"Besök din handelsrådgivare"
"##wage_level_tip##":"Fastställ en lönenivå (ditt folk kommer att jämföra denna med lönerna i Rom)"
"##wages##":"Löner"
"##wait_for_fishing_boat##":"Vi vänta för närvarande på att ett varv skall bygga oss en fiskebåt."
"##waiting_for_free_dock##":"Har kastat ankar, i väntan på ledig kajplats"
"##wall_info##":"Murar skyddar värnlösa medborgare från barbarer. De kan bara motstå en viss grad av attacker, och tjockare murar klarar sig längre."
"##wall##":"Mur"
"##walls_need_a_gatehouse##":"Murar behöver grindstugor, så att vandringsmän och handelsmän kan komma och gå som de vill."
"##warehouse_devastation_mode_text##":"Försöker sända gods till annan plats"
"##warehouse_full_warning##":"VARNING Denna lagerbyggnad är helt fylld. Den kan inte ta emot fler varor."
"##warehouse_gettinfull_warning##":"VARNING Denna lagerbyggnad håller på att bli full. Den kan bara ta emot varor som redan finns, inga nya varutyper."
"##warehouse_info##":"Varor som produceras för handel kräver magasinering. Karavaner besöker handelsmagasinen för att köpa och sälja varor och handelshamnar får sitt gods från intilliggande magasin."
"##warehouse_low_personal_warning##":"Underbemannad. Kan endast sända iväg varor, ej ta emot varor"
"##warehouse_no_workers##":"Endast minimibemanning. Kommer ej att sända eller ta emot varor"
"##warehouse_orders##":"Instruktioner handelsmagasin"
"##warehouse##":"Handelsmagasin"
"##warehouseman##":"Magasinsman"
"##warehouses##":"Handelsmagasin"
"##warning_amphitheater_access##":"Detta hus har inte passerats av en gladiator på ett tag. Det kommer snart att förlora tillgång till amfiteater"
"##warning_barber_access##":"Om ingen barberare går förbi huset snart, kommer det att förlora sin tillgång till barberare"
"##warning_baths_access##":"Om ingen badhusarbetare passerar snart, kommer detta hus att förlora sin tillgång till badhus"
"##warning_college_access##":"Om ingen lärare passerar huset snart, kommer det att förlora sin tillgång till högskola"
"##warning_colloseum_access##":"Detta hus har inte passerats av en lejontämjare på ett tag. Det kommer snart att förlora tillgång till colosseum"
"##warning_doctor_access##":"Om ingen läkare passerar huset snart, kommer det att förlora sin tillgång till läkarklinik"
"##warning_full##":"Varningar PÅ"
"##warning_hippodrome_access##":"Detta hus har inte passerats av en körsven på ett tag. Det kommer snart att förlora tillgång till hippodrom"
"##warning_hospital_access##":"Om ingen kirurg passerar detta hus snart, kommer det att förlora sin tillgång till sjukhus"
"##warning_library_access##":"Om ingen bibliotekarie passerar huset snart, kommer det att förlora sin tillgång till bibliotek"
"##warning_school_access##":"Om inget skolbarn passerar huset snart, kommer det att förlora sin tillgång till skola"
"##warning_some##":"Varningar AV"
"##warning_theater_access##":"Detta hus har inte passerats av en skådespelare på ett tag. Det kommer snart att förlora tillgången till teater"
"##water_build_tlp##":"Byggnader förknippade med vatten"
"##water_caption##":"H2O"
"##water_info##":"Kan inte forceras, men broar kan byggas på vissa platser. Vatten är en vital handelslänk till resten av imperiet via handelshamnar. Lertag måste byggas nära vatten."
"##water_srvc_fountain_and_well##":"Detta område har tillgång till en reservoar via rörledning och dricksvatten från en brunn eller fontän"
"##water_srvc_reservoir##":"Detta område har tillgång till en reservoar via rörledning, vilket gör att fontäner och badhus fungerar"
"##water_srvc_well##":"Detta område har tillgång till dricksvatten"
"##water_supply##":""
"##we_eat_more_thie_produce##":"Vi äter mer än vi producerar"
"##we_eat_much_then_produce##":"Vi äter mycket mer än vi producerar"
"##we_eat_some_then_produce##":"Vi äter något mer än vi producerar"
"##we_produce_less_than_eat##":"Dina invånare äter mer mat än de producerar"
"##we_produce_more_than_eat##":"Vi producerar något mer än vi äter"
"##we_produce_much_than_eat##":"Vi producerar mycket mer än vi äter"
"##we_produce_some_than_eat##":"Vi producerar lagom för att livnära alla"
"##weapon##":"Vapen"
"##weapons_workshop_bad_work##":"Med så få anställda står produktionen nästan still. Det kommer inte att produceras många vapen under det kommande året."
"##weapons_workshop_full_work##":"Denna smedja har alla anställda den behöver, den arbetar fullt ut med att producera vapen."
"##weapons_workshop_info##":"Vapensmeder förvandlar järn till vapen och rustningar, som du kan handla med och göra vinst eller använda för att utrusta dina egna legioner."
"##weapons_workshop_need_resource##":"Denna smedja kräver leverans av järn, från ett magasin eller från ett malmbrott, för att producera vapen."
"##weapons_workshop_need_some_workers##":"Denna smedja är underbemannad, och det tar längre tid att producera vapen än vad det borde."
"##weapons_workshop_no_workers##":"Detta snickeri har inga anställda. Produktionen har upphört."
"##weapons_workshop_patrly_workers##":"Denna smedja utnyttjas inte till maximal kapacitet. Vapenproduktionen kommer att gå något långsammare än vad den borde."
"##weapons_workshop_slow_work##":"Mycket få människor arbetar i smedjan. Som resultat är vapenproduktionen långsam."
"##weapons_workshop##":"Vapensmedja"
"##well_haveno_houses_inarea##":"Denna brunn är överflödig för tillfället, eftersom det inte finns några hus inom dess serviceområde."
"##well_info##":"Medborgare utan tillgång till fontän kan ta vatten från brunnar, men stadsdelar med brunnsvatten är inga trevliga platser att bo på."
"##well##":"Brunn"
"##wharf_full_work##":"Med fullt antal anställda lassar och lossar vi med maximal hastighet."
"##wharf_info##":"Båtar avseglar från fartygsvarvet och hämtar sina besättningar här. Varje fiskehamn kan betjäna en fiskebåt."
"##wharf_our_boat_fishing##":"Vår fiskebåt befinner sig vid fiskevattnet och fångar just nu fisk."
"##wharf_our_boat_return##":"Vår båt seglar mot hamn."
"##wharf_out_boat_ready_fishing##":"Vår fiskebåt seglar ut till fiskevattnen."
"##wharf_out_boat_return_with_fish##":"Vår fiskebåt seglar tillbaka från fiskevattnen med sin fångst."
"##wharf##":"Fiskehamn"
"##wheat_farm_bad_work##":"Det finns mycket få jordbruksarbetare här. Som resultat är veteproduktionen långsam."
"##wheat_farm_full_work##":"Denna lantgård har alla anställda det behöver. Den får maximum avkastning på sin areal."
"##wheat_farm_info##":"Vetekorn är det grundläggande livsmedlet för ditt folk. Det måste lagras i sädesmagasin för att livnära ditt folk, eller i handelsmagasin för export."
"##wheat_farm_need_some_workers##":"Denna lantgård är underbemannad. Arbetarna kan inte så alla de fält som finns."
"##wheat_farm_no_workers##":"Denna lantgård har inga anställda. Jorden ligger i träda."
"##wheat_farm_patrly_workers##":"Denna lantgård arbetar under sin maximala kapacitet. Fler arbetare skulle öka produktiviteten."
"##wheat_farm##":"Veteodling"
"##wheat##":"Vete"
"##win_syracusae_text##":"Bäste ståthållare, det var en lysande uppvisning. Du övertygade grekerna att överge sina planer för Syracusae vilket lägger hela Medelhavet för Roms fötter. Efter en sådan imponerande bragd kommer du aktivt att delta i framtida planer."
"##wine_workshop_bad_work##":"Med så få anställda står produktionen nästan still. Det kommer att produceras mycket lite vin under det kommande året."
"##wine_workshop_full_work##":"Denna vingård har alla anställda den behöver och arbetar fullt ut med att producera vin."
"##wine_workshop_info##":"Vinhandlare förvandlar druvor till vin, vilket patricierna kräver om de skall bygga villor. Vin är en handelsvara som är begärlig för många."
"##wine_workshop_need_resource##":"Denna vingård kan inte producera vin förrän den får en leverans av druvor från ett magasin eller en druvodling."
"##wine_workshop_no_workers##":"Denna vingård har inga anställda. Produktionen har upphört."
"##wine_workshop_slow_work##":"Mycket få människor arbetar vid denna vingård. Som resultat är vinproduktionen långsam."
"##wine_workshop##":"Vingård"
"##wine_workshops_need_some_workers##":"Denna vingård är underbemannad och det tar mycket längre tid att producera vin än vad det borde."
"##wine_workshops_patrly_workers##":"Denna vingård utnyttjar inte full kapacitet. Vinproduktionen något långsammare än vad den borde vara."
"##wine##":"Vin"
"##wnd_ratings_title##":"Ställning"
"##wndrt_culture##":"Kultur"
"##wndrt_favor_tooltip##":"Klicka här för information om din popularitetsställning"
"##wndrt_favour##":"Popularitet"
"##wndrt_need##":"Behövs"
"##wndrt_peace_tooltip##":"Klicka här för information om din fredsställning"
"##wndrt_peace##":"Fredsställning"
"##wndrt_prosperity_tooltip##":"Klicka här för information om din välståndsställning"
"##wndrt_prosperity##":"Välstånd"
"##work##":"I bruk"
"##workers_yearly_wages_is##":"Beräknad årlig kostnad för"
"##working_build_poor_labor_warning##":"Varning: Dålig tillgång till arbetskraft"
"##working_building_need_road##":"VARNING. Denna byggnad fungerar ej. Den ligger inte intill en väg, och dess anställda kommer ej fram"
"##working_have_awesome_labor_access##":"Denna byggnad har för närvarande utmärkt tillgång till arbetskraft"
"##working_have_bad_labor_access##":"Denna byggnad har för närvarande dålig tillgång till arbetskraft"
"##working_have_good_labor_access##":"Denna byggnad har för närvarande god tillgång till arbetskraft"
"##working_have_no_labor_access##":"Denna byggnad har för närvarande ingen tillgång till arbetskraft"
"##working_have_some_labor_access##":"Denna byggnad har för närvarande viss tillgång till arbetskraft"
"##working_have_very_little_labor_access##":"Denna byggnad har för närvarande mycket liten tillgång till arbetskraft"
"##wrath_of_neptune_title##":"Neptuns Vrede"
"##wt_cartPusher##":"Vagndragare"
"##wt_criminal##":"Brottsling"
"##wt_emigrant##":""
"##wt_endeavor##":"Endeavor"
"##wt_engineer##":""
"##wt_gladiator##":"Gladiator"
"##wt_homeless##":"Hemlös"
"##wt_immigrant##":"Immigrant"
"##wt_indigene##":"Inföding"
"##wt_legioanry##":"Legionär"
"##wt_librarian##":"Bibliotekarie"
"##wt_lion_tamer##":"Lejontämjare"
"##wt_marketBuyer##":"Marknadsbesökare"
"##wt_marketLady##":"Marknadshandlare"
"##wt_missionary##":"Missionär"
"##wt_missioner_average_life##":"Var hälsad! Jag ser att det finns mycket att göra med att lära dessa barbarer fördelarna med Roms välvilja."
"##wt_missioner_normal_life##":"Jag är så glad att vara romare. Du skulle se vad dessa barbarer håller på med i sina hyddor!"
"##wt_prefect##":"Prefekt"
"##wt_priest##":"Präst"
"##wt_rioter##":"Upprorsman"
"##wt_sheep##":"Får"
"##wt_surgeon##":"Kirurg"
"##wt_taxCollector##":"Skatteindrivare"
"##wt_teacher##":"Lärare"
"##wt_wolf##":"Varg"
"##year##":"Sädesmagasin lagrar"
"##years##":"Sädesmagasin lagrar"
"##yes##":"Ja"
"##your_favor_is_dropping_catch_it##":"Din popularitet i Rom minskar. Du måste fånga Caesars intresse på ett eller annat sätt!"
"##your_favour_increased_from_last_year##":"Din ställning i Rom har förbättrats sedan förra året."
"##your_favour_unchanged_from_last_year##":"Din ställning är oförändrad sedan förra året."
"##your_prosperity_raising##":"Din välståndsställning förbättras."
"##your_province_quiet_and_secure##":"Din provins lugna och säkra tillvaro har blivit legendarisk. Andra ståthållare planerar förmodligen att dra sig tillbaka hit!"
"##your_salary_frowned_senate##":"I Rom ser man ner på din fräckhet att betala dig själv en lön som är högre än din rang."
"#winning_population##":"Vinnande befolkning"
"Variable":"SVENSKA (v1.0)"










































































































































































































































































































































































































































}
