{
"##some_food_on_next_month##":"- vissa livsmedel till kommande månad"
"##have_no_food_on_next_month##":"- inga livsmedel till kommande månad"
"##dn_for_open_trade##":"för att öppna handelsväg"
"##small_food_on_next_month##":"- mycket lite mat till kommande månad"
"##no_target_population##":"( Ingen målbefolkning )"
"##teacher_good_life##":"Staden får full pott. Det är en underbar plats."
"##actor_gods_angry##":"Aaagh!! Gudarna är rasande. Vi går under!"
"##ovrm_academy##":"Högskola"
"##academy##":"Högskola"
"##accept##":"Acceptera"
"##accept_goods##":"Acceptera varor"
"##accept_promotion##":"Acceptera befordran"
"##accept_deity_status##":"Acceptera ställningen som kejsare!"
"##accepting##":"Accepterar"
"##bath_access##":"Badtillgång"
"##barber_access##":"Barberartillgång"
"##academy_full_work##":"Denna högskola används, och ungdomarna i stadsdelen lär sig sociala färdigheter."
"##aqueduct_no_water##":"Denna akvedukt transporterar inte vatten mellan reservoarer eftersom den saknar vattenkälla."
"##also_fountain_in_well_area##":"Denna brunn är överflödig för tillfället, eftersom alla hus som den betjänar tar sitt vatten från en fontän."
"##academy_no_workers##":"Denna högskola används inte, och är därför värdelös för lokalsamhället."
"##baths_need_reservoir##":"Detta badhus behöver en rörledning till en reservoar."
"##baths_full_work##":"Detta badhus används, besökarna blir rena och avslappnade."
"##baths_no_workers##":"Detta badhus används inte, och är därför värdelöst för lokalsamhället."
"##avesome_library_access##":"Detta hus har nyligen passerats av en bibliotekarie. Det kommer att ha tillgång till bibliotek under lång tid framåt"
"##avesome_hospital_access##":"Detta hus passerades nyligen av en kirurg. Det kommer att ha tillgång till sjukhus under lång tid framåt"
"##avesome_amphitheater_access##":"Detta hus passerades nyligen av en gladiator. Det kommer att ha tillgång till amfiteater under lång tid framåt"
"##avesome_colloseum_access##":"Detta hus passerades nyligen av en lejontämjare. Det kommer att ha tillgång till ett colosseum under lång tid framåt"
"##avesome_clinic_access##":"Detta hus passerades nyligen av en läkare. Det kommer att ha tillgång till en klinik under lång tid framåt"
"##avesome_college_access##":"Detta hus passerades nyligen av en lärare. Det kommer att ha tillgång till högskola under lång tid framåt"
"##avesome_hippodrome_access##":"Detta hus har nyligen passerats av en körsven. Det kommer att ha tillgång till hippodrom under lång tid framåt"
"##bath_no_access##":"Detta hus har inte tillgång till ett fungerande badhus"
"##amphitheater_no_access##":"Detta hus har inte tillgång till en amfiteater"
"##building_need_road_access##":"Denna byggnad behöver tillgång till väg"
"##actorColony_no_workers##":"Denna koloni är övergiven. Utan tillgång till mentorer kan inga nya skådespelare utbildas."
"##0_entertainment_access##":"Denna boning har inte tillgång till underhållning överhuvudtaget"
"##clay_pit_full_work##":"Detta lertag har alla anställda det behöver, och arbetar fullt ut med att producera lera."
"##clay_pit_need_some_workers##":"Detta lertag utnyttjar inte full kapacitet. Som resultat kommer lerproduktionen att gå något långsammare."
"##clay_pit_no_workers##":"Detta lertag har inga anställda. Produktionen har upphört."
"##clay_pit_patrly_workers##":"Detta brott är underbemannat, och det tar längre tid än det borde att producera marmorn."
"##avesome_theater_access##":"Detta hus passerades nyligen av en skådespelare. Det kommer att ha tillgång till teater under lång tid framåt"
"##awesome_baths_access##":"Detta hus har tillgång till badhus"
"##awesome_barber_access##":"Detta hus har tillgång till barberare"
"##avesome_school_access##":"Detta hus passerades nyligen av ett skolbarn. Det kommer att ha tillgång till skola under lång tid framåt"
"##amphitheater_no_workers##":"Denna amfiteater är stängd. Den har inga anställda, och erbjuder ingen förströelse åt det lokala samhället."
"##amphitheater_have_only_battles##":"Denna amfiteater erbjuder gladiatorkamp som förströelse. Den söker skådespelare för att sätta upp några pjäser."
"##amphitheater_have_never_show##":"Denna amfiteater har sällan några föreställningar. Den behöver skådespelare och gladiatorer."
"##amphitheater_full_work##":"Denna amfiteater erbjuder sitt samhälle både intressant gladiatorkamp och pjäser med lokala skådespelare."
"##amphitheater_have_only_shows##":"Denna amfiteater sätter upp pjäser med lokala aktörer. Den kan attrahera större publik om den även har gladiatorer."
"##aqueduct_work##":"Denna akvedukt transporterar vatten mellan reservoarer."
"##citizen_gods_angry3##":"Den här ståthållaren har ingen respekt för gudarna."
"##engineer_need_workers##":"Staden skulle fungera bättre om det fanns nog med arbetare."
"##citizen_need_workers5##":"Staden behöver fler arbetare!"
"##romeGuard_need_workers##":"Den här staden behöver många fler arbetare."
"##taxCollector_need_workers##":"Den här staden behöver fler arbetare och det genast."
"##citizen_need_workers3##":"Staden lider stor brist på arbetare."
"##priest_need_workers##":"Detta ställe behöver många fler arbetare."
"##scholar_low_entertainment##":"Staden är så tråkig. Jag vill se fler föreställningar."
"##barber_no_access##":"Detta hus har inte tillgång till en barberare"
"##citizen_gods_angry##":"Detta är en hednisk stad. Den behöver fler tempel."
"##marketBuyer_low_entertainment##":"Detta måste vara den tråkigaste staden i imperiet."
"##actor##":"Skådespelare"
"##administration_building##":"Administrativa- eller regeringsbyggnader"
"##mainmenu_package##":"Advancerade inställningar"
"##package_options##":"Avancerade inställningar"
"##month_8_short##":"Ago"
"##advemployer_panel_title##":"Arbetstilldelning"
"##immigrant_want_to_be_liontamer##":"Jag har hört att det finns arbete här. Jag vill bli lejontämjare."
"##amphitheatres##":"Amfiteatrar"
"##ovrm_amphitheater##":"Amfiteatrar"
"##amphitheater##":"Amfiteater"
"##adve_entertainment##":"Underhållning"
"##entertainment_advisor_title##":"Underhållning"
"##bathlady##":"Badarbetare"
"##barracks_need_some_workers##":"Pga. personalbrist utbildar vi nya soldater långsammare än vanligt men vi har de vapen som krävs för att utbilda alla typer av soldater."
"##barracks_full_work##":"Vi utbildar nya soldater med maximal effektivitet och vi har vapen för att utbilda alla typer av soldater."
"##cancel##":"Avbryt"
"##cancelBtnTooltip##":"Avbryt denna operation"
"##aqueduct##":"Akvedukt"
"##aqueduct_info##":"Akvedukter gör det möjligt att konstruera reservoarer långt från vatten, vilket gör det möjligt för fontäner att förse staden med vatten."
"##month_4_short##":"Apr"
"##cartPusher_cantfind_destination##":"Det skulle gå snabbare att dra varorna till Rom än dit jag ska."
"##arrange_festiable_for_this_god##":"Arrangera en festival till denna guds ära"
"##btn_showprice_tooltip##":"Visar import-/exportpriser för alla varor, som anbefallt av Rom"
"##city_need_workers_title##":"Behöver fler arbetare"
"##clay##":"Lera"
"##clay_pit_info##":"Tag lera och handla med, eller leverera den till krukmakerier. Folket behöver krukor för att bebo Insulaen."
"##clay_factory_stock##":"Lagrad lera,"
"##architect##":"Arkitekt"
"##arabian_stallions##":"Arabiska hingstar"
"##advchief_military##":"Militär"
"##adve_military##":"Militär"
"##mainmenu_dlc_articles##":"Artiklar"
"##barbarian_attack_title##":"Barbarer anfaller!"
"##clay_pit_bad_work##":"Med nästan inga grävare vid detta lertag, står produktionen nästan helt still. Det kommer inte att produceras mycket lera under det kommande året."
"##having_some_slums_lack_migration##":"Att ha slumområden förhindrar immigration"
"##actorColony_patrly_workers##":"Vi har bara halva personalstyrkan, och kan därför endast utbilda en skådespelare under nästa månad."
"##charioteer_school_patrly_workers##":"Vi har bara halva personalstyrkan, och kan därför endast tillverka en vagn under nästa månad."
"##actorColony_slow_work##":"Vi lider av svår personalbrist, och kommer att få kämpa för att utbilda en ny skådespelare under de kommande två månaderna."
"##chatioteer_school_slow_work##":"Vi lider av svår personalbrist, och kommer att få kämpa för att bygga en enda ny vagn under de kommande två månaderna."
"##ovrm_baths##":"Bad"
"##baths##":"Badhus"
"##bath_1##":"Badhus"
"##bath##":"Badhus"
"##balance##":"Balans"
"##ballista##":"Katapult"
"##barracks##":"Förläggningar"
"##wn_barbarian##":"Barbar"
"##ovrm_barber##":"Barberare"
"##wharf_info##":"Båtar avseglar från fartygsvarvet och hämtar sina besättningar här. Varje fiskehamn kan betjäna en fiskebåt."
"##britons##":"Britter"
"##mediolanum_win_text##":"Att Hannibal kunde korsa Alperna med sina elefanter var häpnadsväckande. Att Mediolanum skulle blomstra trots hans attacker är ett mirakel. Din framgång vände lyckan i det puniska kriget till Roms fördel. Hela Rom tackar dig."
"##caesar_assign_new_title##":"Caesar har befordrat dig till graden"
"##native_field##":"Ängmark"
"##big_hut##":"Stort hus"
"##patrician_high_workless##":"Detta är skandalöst. Jag har aldrig sett så många arbetslösa plebejer."
"##ceres_goodmood_info##":"Ceres skänker fruktsamhet åt jorden, och får plantorna att växa. Blidka henne, eller bered dig på hungersnöd."
"##patrician_low_entertainment##":"Medborgare! Är icke detta den tråkigaste staden i riket?"
"##citizen_are_rioting##":"Medborgarna gör uppror!"
"##quaestor##":"Kvestor"
"##city_cyrene##":"Cyrene"
"##advice_at_culture##":"Klicka här för information om din kulturställning"
"##taxСollector_low_tax_collected##":"Att driva in skatt från dessa hårt arbetande människor får mig nästan att gråta - men bara nästan!"
"##actorColony##":"Skådespelarkoloni"
"##advpopulation_text_census##":"Befolkningssammansättning efter ålder (år)"
"##advpopulation_text_society##":"Befolkningssammansättning efter inkomst"
"##fired##":"Avskedad!"
"##mainmenu_dlc_concepts##":"Begrepp"
"##animal_contests_run##":"Djurtävlingarna pågår ytterligare"
"##chief_advisor##":"Huvudrådgivare"
"##advisors##":"Senat"
"##buildings##":"Byggnation"
"##build_road_tlp##":"Bygg vägar"
"##build_housing##":"Bygg bostäder"
"##clay_pit_need_close_to_water##":"Bygg lertag nära vattnet"
"##build_markets_to_distribute_food##":"Bygg marknader för att distribuera maten som lagrats här"
"##build_fishing_boat##":"Vi bygger båtar på beställning från en fiskehamn i staden."
"##children##":"Barn"
"##school_info##":"Barn måste gå i stadsdelsskolorna för att lära sig grunderna i läsning, skrivning och retorik om de skall kunna växa upp till produktiva vuxna."
"##big_tent##":"Stort tält"
"##mainmenu_credits##":"Credits"
"##engineering_post_no_workers##":"Utan egna anställda ingenjörer, denna byggnad  riskerar att falla samman."
"##militaryAcademy_no_workers##":"Utan personal kan vi inte finslipa kunskaperna för stadens nya soldater. De tvingas att gå direkt till sina poster och hoppas på det bästa."
"##fort_legionaries_no_workers##":"Utan personal kan vi inte utbilda en enda ny rekryt. Mars hjälpe oss i krigstid!"
"##marketBuyer_high_workless##":"Med denna höga arbetslöshet måste jag arbeta hårt för att behålla mitt jobb."
"##barracks_bad_weapons_bad_workers##":"Med minimal personal och utan vapen i lager, får vi kämpa för att utbilda till och med de mest enkla trupper."
"##ad##":"eKr"
"##age_ad##":"eKr"
"##charioter_so_hungry##":"Hungrig? Jag kan äta en häst, så lite mat finns det."
"##immigrant_so_hungry##":"Om jag stannar längre dör jag. Det finns ingen mat någonstans."
"##citizen_high_workless2##":"Om jag inte får arbete snart, måste jag flytta till en annan stad."
"##doctor_gods_angry##":"Om vi inte respekterar gudarna mer, kommer vi att få känna på deras vrede."
"##city_damascus##":"Damascus"
"##city_have_goods_for_request##":"Dina lager rapporterar att du nu har tillräckligt av dessa varor för att uppfylla begäran från kejsaren."
"##hospital_info##":"Även om ingen vill bo i närheten av dem, räddar sjukhus liv. Staden borde ha tillräckligt med sängplatser för alla sina invånare."
"##cartpusher_cant_unload_goods_in_factory##":"...ta emot dem. Jag har hört att de behöver mer arbetskraft."
"##population_registered_as_taxpayers##":"av befolkningen är skatteskrivna"
"##dn's##":"Avsluta byggare"
"##advemployer_panel_denaries##":"dn"
"##road_paved_caption##":"Stenbelagdväg"
"##barber_need_colloseum##":"Efter en dag med rakning och klippning vill jag se en trevlig lejonstrid. Men det går inte att uppbringa här."
"##engineer_low_entertainment##":"Efter en hård dags arbete vill jag se en bra pjäs eller strid. Det finns inte mycket chans till det i den här staden."
"##aedile##":"Edil"
"##clear_land##":"Röj marken"
"##gladiator_need_workers##":"Det är hemskt. Jag har aldrig sett så många lediga jobb."
"##doctor_need_workers##":"Var hälsad! Det saknas många arbetare här."
"##teacher_need_workers##":"Otroligt att det finns så många arbetstillfällen här."
"##really_destroy_fort##":"Är du säker på att du vill ta detta fort ur aktiv tjänst?"
"##tingis_win_text##":"Är du ståthållare eller general? Din utmärkta insats vid Tingis befriar mina legioner från tjänstgöring i väst och låter mig ägna tiden åt andra strävanden. Du börjar bli en nyckelperson i min planering."
"##workers_yearly_wages_is##":"Beräknad årlig kostnad för"
"##meadow_caption##":"Äng"
"##chatioteer_school_no_workers##":"Utan hantverkare kan inga nya vagnar produceras. Som resultat kan hippodromen, om den är i drift, bli lidande."
"##bldm_farm##":"Jordbruk"
"##gmenu_file##":"Arkiv"
"##file##":"Arkiv"
"##scholar_high_workless##":"Det är jättemånga som söker arbete här."
"##employers##":"Anställd arbetsstyrka"
"##fortification##":"Befästning"
"##barber##":"Barberare"
"##barber_full_work##":"Denna barberarlokal används, och ortsbefolkningen är vältrimmad."
"##barber_no_workers##":"Denna barberarlokal används inte, och är därför värdelös för lokalsamhället."
"##barber_shop##":"Barberarsalong"
"##barbers##":"Barberarsalonger"
"##clerk##":"Bokhållare"
"##angry##":"Arga"
"##granery##":"Sädesmagasin"
"##granary_holds##":"Sädesmagasin innehåller"
"##granaries_holds##":"Sädesmagasiner innehåller"
"##adve_administration_religion##":"Styrelse/Religion"
"##win_syracusae_text##":"Bäste ståthållare, det var en lysande uppvisning. Du övertygade grekerna att överge sina planer för Syracusae vilket lägger hela Medelhavet för Roms fötter. Efter en sådan imponerande bragd kommer du aktivt att delta i framtida planer."
"##age_bc##":"BC"
"##bc##":"fKr"
"##exit##":"Avsluta"
"##quit##":"Avsluta"
"##cartPusher_so_hungry##":"...dagen kräver styrka. Hur ska en vagndragare kunna arbeta utan mat?"
"##advchief_haveprofit##":"Tillgångarna har i år stigit med"
"##advchief_havedeficit##":"Tillgångarna har i år minskat med"
"##damascus_win_text##":"Ännu en gång har du uppnått vad svagare män kallar omöjligt. Hela östern åsåg din balansgång i Damaskus. Nu kan jag tryggt hämta hem några av mina syriska legioner."
"##ovrm_aborigen##":"Aborigin"
"##adve_industry_and_trade##":"Industri och handel"
"##advanced_houseinfo##":"Avancerad information om detta hus"
"##adve_engineers##":"Konstruktion"
"##big_domus##":"Stor Insula"
"##return_2_fort##":"Återvänd till fortet"
"##teacher_average_life##":"Jag ger staden åtta av tio poäng."
"##gmenu_exit_game##":"Avsluta spel"
"##gmenu_file_exit##":"Avsluta spel"
"##mainmenu_quit##":"Avsluta spel"
"##city_need_workers_text##":"Din stad behöver fler arbetare"
"##teacher_low_entertainment##":"Staden är så tråkig! Den behöver mer underhållning."
"##teacher_so_hungry##":"Det saknas livsmedel här. Det gör medborgarna olyckliga."
"##exit_without_saving_question##":"Avsluta utan att spara?"
"##gmenu_file_mainmenu##":"Avsluta till huvudmenyn"
"##exit_this_panel##":"Avsluta denna panel"
"##cartPusher_normal_life##":"Allt verkar fungera bra här."
"##more_person##":"Anställd"
"##more_people##":"Anställda"
"##bldm_factory##":"Verkstäder"
"##army_marker##":"Armémarkör"
"##bldm_raw_material##":"Råmaterial"
"##mainmenu_mcmxcviii##":"MCMXCVIII"
"##clay_pit##":"Lertag"
"##advemployer_panel_haveworkers##":"arbete"
"##abwrk_working##":"fungerar"
"##labor##":"Arbetskraft"
"##actor_low_entertainment##":"Jag arbetar så hårt jag förmår, men underhållningen i staden räcker inte till på långa vägar."
"##advemployer_panel_workers##":"arbetare"
"##actorColony_need_some_workers##":"Vi är något underbemannade, och kan därför endast utbilda två nya skådespelare per månad."
"##charioteer_school_need_some_workers##":"Vi är något underbemannade, och kan därför endast tillverka två nya vagnar per månad."
"##wndrt_need##":"Behövs"
"##ceres_badmood_info##":"Ceres missnöje är farligt, eftersom hon skyddar folket från dåliga skördar och hungersnöd."
"##advemployer_panel_needworkers##":"behöver"
"##requierd##":"Behov"
"##citizen_low_salary##":"Min hund skulle inte arbeta för de löner de betalar här. Jag ger mig av."
"##amphitheater_haveno_gladiator_bouts##":"Ingen gladiatorkamp för närvarande"
"##amphitheater_haveno_shows##":"Inga pjäser för närvarande"
"##barber_info##":"Ingen civiliserad man visar sig orakad offentligt! Alla medborgare behöver regelbundet besöka en barberare för att kunna avancera i samhället."
"##barracks_info##":"Ingen kan gå med i en romersk legion utan att först komma hit. Alla nya rekryter kommer hit."
"##citizen_good_education##":"Den här staden är mer kultiverad än någon annan i riket!"
"##abwrk_not_working##":"fungerar inte"
"##citizen_low_entertainment4##":"Man kan inte roa sig alls på det här stället!"
"##citizen_high_workless4##":"Jag har aldrig sett så många arbetslösa medborgare förut."
"##actorColony_bad_work##":"Jag har ingen personal utöver mig själv. Jag kan inte arbeta under dessa förhållanden! Som bäst kan jag utbilda en skådespelare på tre månader."
"##chatioteer_school_bad_work##":"Jag har ingen personal utöver mig själv. Jag kan inte arbeta under dessa förhållanden! Jag kan bara bygga en vagn på tre månader."
"##prefect_high_workless##":"Jag har aldrig sett så många arbetslösa!"
"##advlegion_norequest##":"Vi har inte fått någon begäran om hjälp från imperiet"
"##advlegion_noalarm##":"Vi har inga rapporter om hot mot staden"
"##barber_average_life##":"Är inte den här staden ett riktigt klipp?"
"##cartPusher_low_entertainment##":"...vagnar. Det är mer underhållande än resten av den här staden."
"##cant_demolish_bridge_with_people##":"Kan inte förstöra bro med människor på"
"##cartPusher_gods_angry##":"...religiös, men inte ens jag skulle behandla gudarna på det här sättet."
"##barber_so_hungry##":"En hårklippning får dig att glömma hungern. Och det är många hungriga i den här staden."
"##baths_info##":"Civiliserade människor badar minst en gång om dagen. Utöver bättre hälsa utgör baden även en önskvärd träffpunkt med olika rekreativa aktiviteter."
"##advchief_employment##":"Arbete"
"##gmenu_options##":"Alternativ"
"##mainmenu_options##":"Alternativ"
"##city##":"Stad"
"##city_need_more_workers##":"Din stad kräver fler arbetare"
"##city_has_debt##":"Staden har en skuld till Rom på"
"##empmap_distant_romecity_tip##":"Avlägsen romersk stad"
"##city_has_runout_debt##":"Din stad har inga pengar kvar. Caesar har gått med på att ge dig mer, men han kommer inte vara så generös nästa gång. Exportera varor för att generera mer inkomst till din stad."
"##big_palace##":"Stort palats"
"##target_population_is##":"( Målbefolkningen är"
"##prosperity_lack_that_you_pay_less_rome##":"Att betala lägre löner än Rom ger din stad rykte att vara mindre blomstrande."
"##gladiator_low_entertainment##":"Tråkigt! Det säger alla om det här stället, trots mina tappra insatser. Staden behöver verkligen mer underhållning."
"##bridge##":"Bro"
"##bridges##":"Broar"
"##population_tooltip##":"Befolkningsmängd"
"##mission_wnd_population##":"Befolkning"
"##population##":"Befolkning"
"##advpopulation_title_population##":"Befolkning - Historia"
"##advpopulation_title_census##":"Befolkning - Folkräkning"
"##advpopulation_title_society##":"Befolkning - Samhälle"
"##adve_prefectures##":"Prefekturer"
"##advemployer_panel_priority##":"prioritering"
"##adve_food##":"Livsmedelsproduktion"
"##chatioteer_school##":"Skola för körsvenner"
"##chatiotSchool##":"Skola för körsvenner"
"##bolt##":"Armborst"
"##actor_so_hungry##":"Jag kan inte uppträda utan mer mat."
"##tower_may_build_on_thick_walls##":"Du kan endast bygga torn på tjocka murar"
"##access_ramp##":"Åtkomstramp"
"##reorient_map_to_north##":"Ändra visningen norrut"
"##reject##":"Avvisa varor"
"##return_to_main_map##":"Återvänd till spelets huvudkarta"
"##advemployer_panel_romepay##":"Rom betalar"
"##arrow##":"Pil"
"##architect_salary##":"Arkitektlön på"
"##caesar_salary##":"Caesars lön på"
"##citizen_salary##":"Medborgarlön på"
"##clerk_salary##":"Bokhållarlön på"
"##adve_health_education##":"Hälsa och utbildning"
"##mainmenu_plname##":"Ändra namn"
"##increase_trading_title##":"Begär ändringar"
"##edadv_need_better_access_school_or_colege##":"Bättre skola eller högskola och tillgång till bibliotek skulle förbättra vissa områden i staden. Man skall inte behöva gå långt för att lära sig något!"
"##advemployer_panel_sector##":"Sektor"
"##adve_water##":"Vattenförsörjning"
"##senatepp_unemployment##":"Arbetslöshet"
"##advemployer_panel_workless##":"Arbetslös arbetsstyrka "
"##citizen_high_workless10##":"Arbetslösheten är så hög att hela staden mår dåligt."
"##cartPusher_high_workless##":"...min fru har slutat tjata om att jag ska skaffa mig ett nytt arbete."
"##barber_high_workless##":"Arbetslösheten är så hög att den får håret att stå på ända!"
"##doctor_high_workless##":"Arbetslösheten är mycket hög. Jag funderar på att ge mig av."
"##actor_high_workless##":"Det är så stor arbetslöshet att jag inte förmår lära mig mina repliker."
"##priest_high_workless##":"Arbetslösheten är oroväckande hög"
"##migration_lack_workless##":"Arbetslöshet minskar antalet immigranter."
"##citizens_additional_rooms_for##":"Extra utrymme för"
"##teacher_high_workless##":"Bara jag inte förlorar jobbet. Arbetslösheten är så hög att jag inte skulle få ett nytt."
"##send_legion_to_emperor##":"Be din militära rådgivare att avdela några stridsklara legioner i imperiets tjänst"
"##adjust_tax_rate##":"Justera skattenivån i staden"
"##adjust_exact##":"Ställ in den exakta summa du vill donera"
"##city_health##":"Hälsosituation"
"##advlegion_window_title##":"Legionstatus"
"##advchief_food_stocks##":"Matförråd"
"##academy_trained##":"Utbildad på högskola"
"##below_average##":"Under medel"
"##scrw_subject##":"Ämne"
"##city_sounds_on##":"Stadsljud är på"
"##city_sounds_off##":"Stadsljud är av"
"##scholar_so_hungry##":"Jag svälter ihjäl!"
"##engineer_high_workless##":"Jag har tur som har ett arbete i denna tid av arbetslöshet."
"##recruter_gods_angry7##":"Vi har problem! Gudarna är förargade på oss."
"##priest_gods_angry##":"Vi är i fara! Staden visar ingen respekt för gudarna."
"##actorColony_full_work##":"Det är med nöje vi tillkännager att vi, med full sysselsättning, kan hjälpa upp till fyra nya skådespelare varje månad."
"##charioteer_school_full_work##":"Det är med nöje vi tillkännager att vi, med full sysselsättning, kan slutföra upp till fyra nya vagnar varje månad."
"##mainmenu_dlc_wallpapers##":"Bakgrundsbilder"
"##clear_land_caption##":"Tomt land"
"##hold_ceres_festival##":"Anordna festival för Ceres"
"##hold_mars_festival##":"Anordna festival för Mars"
"##hold_mercury_festival##":"Anordna festival för Merkurius"
"##hold_neptune_festival##":"Anordna festival för Neptunus"
"##hold_venus_festival##":"Anordna festival för Venus"
"##new_festival##":"Anordna ny festival"
"##education_awesome##":"Alla som kräver utbildningsmöjligheter i staden har dem, och dessa är perfekta i hela staden."
"##doctor_so_hungry##":"Folk är undernärda, men det saknas mat att bota det med."
"##ovrm_education##":"Allt"
"##ovrm_entrertainment##":"Allt"
"##colege_access_perfectly##":"Alla områden som kräver utbildningsmöjligheter har tillgång till dem, men fler högskolor skulle minska storleken på klasserna."
"##library_access_perfectrly##":"Alla områden som kräver utbildningsmöjligheter har tillgång till dem, men fler bibliotek skulle minska trängseln."
"##school_access_perfectly##":"Alla områden som kräver utbildningsmöjligheter har tillgång till dem, men fler skolor skulle minska storleken på klasserna."
"##romeGuard_average_life##":"Allt verkar lugnt här."
"##engineer_average_life##":"Allt tycks fungera väl här."
"##become_trade_center##":"Utse till handelscentral"
"##city_have##":"Stadens skattkammare har tillgångar på"
"##tower##":"Torn"
"##age_uc##":"UC"
"##seamrchant_another_successful_voyage##":"Ännu en lyckosam resa. Förtjänsten från denna stad gör att man står ut med sjösjukan."
"##briton##":"En britt"
"##egift_chest_of_sapphire##":"En kista med safirer"
"##captured_city##":"En erövrad stad"
"##barber_good_life##":"Rakning eller klippning, medborgare? Livet här är lätt att leva, inte sant?"
"##barbarian_warrior##":"En barbarisk soldat"
"##carthaginian_soldier##":"En karthagisk soldat"
"##road_paved_title##":"En finare typ av väg"
"##use_and_trade_resource##":"Använder och byteshandlar med denna vara"
"##actor_average_life##":"Livet här är helt enkelt ljuvligt."
"##priest_good_life##":"Livet är mycket behagligt i denna stad."
"##big_villa##":"Stor villa"
"##charioteer##":"Körsven"
"##teacher_gods_angry##":"Vi får känna gudarnas vrede om vi inte bygger fler tempel snart."
"##engineer_gods_angry##":"Måtte gudarna vara mig nådiga. Det är inte mitt fel att ståthållaren hånar dem."
"##romeGuard_gods_angry##":"Gudarna är rasande över denna plats!"
"##barber_gods_angry##":"Gudarna är rasande. Jag önskar att ståthållaren kunde bygga fler tempel."
"##wt_romeHorseman##":"Beridna stödtrupper"
"##visit_labor_advisor##":"Besök din arbetsrådgivare"
"##visit_population_advisor##":"Besök din befolkningsrådgivare"
"##visit_financial_advisor##":"Besök din finansrådgivare"
"##visit_health_advisor##":"Besök din hälsorådgivare"
"##visit_trade_advisor##":"Besök din handelsrådgivare"
"##visit_chief_advisor##":"Besök din huvudrådgivare"
"##visit_imperial_advisor##":"Besök din imperierådgivare"
"##visit_military_advisor##":"Besök din militärrådgivare"
"##visit_religion_advisor##":"Besök din religionsrådgivare"
"##visit_rating_advisor##":"Besök din ställningsrådgivare"
"##visit_entertainment_advisor##":"Besök din underhållningsrådgivare"
"##visit_education_advisor##":"Besök din utbildningsrådgivare"
"##pay_to_open_trade_route?##":"Betala för att öppna denna väg?"
"##emp_pay_open_this_route_question##":"Betala för att öppna denna väg?"
"##library##":"Bibliotek"
"##libraries##":"Bibliotek"
"##ovrm_library##":"Bibliotek"
"##wt_librarian##":"Bibliotekarie"
"##mainmenu_video##":"Bildskärmsinställningar"
"##screen_settings##":"Bildskärmsinställningar"
"##blood_sports_add_spice_to_life##":"Blodsporter ger krydda åt alla."
"##egift_modest##":"Blygsam:"
"##replay_game##":"Börja om denna karta"
"##devastate_warehouse##":"BÖRJA tömma magasin"
"##god_good##":"Bra"
"##lumber_mill##":"Brädgård"
"##ovrm_fire##":"Brand"
"##fire##":"Brand"
"##burning_ruins##":"Brinnande ruin"
"##migration_people_away##":"Brist på arbete driver bort människor"
"##migration_middle_lack_workless##":"Hög arbetslöshet är ett problem"
"##migration_lack_empty_house##":"Brist på husrum begränsar immigrationen"
"##migration_lessfood_granary##":"Brist på livsmedel i sädesmagasinen minskar immigrationen"
"##migration_empty_granary##":"Brist på mat förhindrar immigration"
"##migration_low_food_stocks##":"Bristen på mat är ett problem"
"##ovrm_crime##":"Brott"
"##advchief_crime##":"Brott"
"##layer_crime##":"Brott"
"##low_crime_risk##":"Brott inträffar sällan i detta område"
"##advchief_which_crime##":"Brottsligheten håller på att bli ett problem."
"##wt_criminal##":"Brottsling"
"##prefect_low_entertainment##":"Brottslingarna jag tar får bättre underhållning än den här staden!"
"##well##":"Brunn"
"##iron_mine_info##":"Bryt järn för att handla med, eller för att leverera till vapensmedjorna. Utrusta din armé med hemgjorda vapen, eller exportera dem till andra provinser."
"##quarry_info##":"Bryt marmor ur intilliggande klippor och använd den till att bygga orakel och stora tempel. Marmor är vanligen en värdefull exportvara."
"##timber_mill_need_trees##":"Bygg brädgård intill träden"
"##need_timber_mill##":"Bygg en brädgård"
"##colloseum_haveno_gladiatorpit##":"Bygg en gladiatorskola för att arrangera matcher här"
"##need_iron_mine##":"Bygg en järngruva"
"##need_olive_farm##":"Bygg en olivodling"
"##need_actor_colony##":"Bygg en skådespelarkoloni för att sända skådespelare hit"
"##need_charioter_school##":"Bygg en skola för körsvenner för att se kapplöpningar"
"##need_vines_farm##":"Bygg en vingård"
"##need_lionnursery##":"Bygg ett lejonhus för att arrangera djurtävlingar"
"##farm_need_farmland##":"Bygg jordbruk på jordbruksmark (leta efter gult gräs)"
"##build_senate_for_advisors##":"Bygg senatorbyggnad"
"##ovrm_build##":"Byggnad"
"##health_advisor##":"Byggnader förknippade med hälsa"
"##water_build_tlp##":"Byggnader förknippade med vatten"
"##emperor_changed_title##":"Byte av kejsare"
"##сaesar##":"Caesar"
"##emperoradv_caesar_has_high_respect_for_you##":"Caesar respekterar dig mer än någon annan ståthållare någonsin!"
"##capua_title##":"Capoue: une province pacifique"
"##carthago_title##":"Carthago: une province dangereuse"
"##god_ceres_short##":"Ceres"
"##smallcurse_of_ceres_description##":"Ceres är missnöjd med din brist på vördnad och ödelägger hela din skörd som en varning till dig."
"##smallcurse_of_ceres_title##":"Ceres är upprörd"
"##wrath_of_ceres_title##":"Ceres vrede"
"##small_ceres_temple##":"Cerestempel"
"##caesarea_title##":"Césarée: province équitablement pacifique"
"##god_charmed##":"Charmerade"
"##ovrm_colloseum##":"Colleseum"
"##colloseum##":"Colosseum"
"##colloseums##":"Colosseum"
"##colloseum_info##":"Colosseum och amfiteatrar behöver alltid nya gladiatorer för att ersätta förlorarna."
"##corinthus##":"Corinthus"
"##day##":"Dag"
"##days##":"Dagar"
"##god_poor##":"Dålig"
"##poor_housing_discourages_migration##":"Dåliga bostäder motverkar invandring trots välståndet i staden"
"##city_fire_text##":"Dåligt underhåll har gjort att det börjat brinna. Just nu sveper elden genom olika områden i staden."
"##damascus_title##":"Damaskus: en relativt farlig provins"
"##date_tooltip##":"Datum"
"##date##":"Datum"
"##scrw_date##":"Datum"
"##gladiator_high_workless##":"De arbetslösa är så många här. Jag önskar vi kunde få träna oss på några av dem."
"##house_not_report_about_crimes##":"De boende har inte rapporterat någon brottslighet."
"##greatPalace_info##":"De boende i detta palats befinner sig högst upp i det romerska samhället. De saknar inte något. Bara att lyckas hålla dem nöjda är en storartad insats."
"##chatioteer_school_info##":"De hantverkare som arbetar här bygger snabba, kraftiga vagnar och utbildar förarna. Kapplöpningarna i hippodromen är mycket populära."
"##city_under_rome_attack##":"De legioner från imperiet som närmar sig skrämmer dina invånare och förbättrar inte din fredsställning."
"##immigrant_much_food_here##":"De påstår att det finns mat här. Är det en bra plats att bo på?"
"##month_12_short##":"Dec"
"##wt_rprotestor##":"Demonstrant"
"##scholar_good_life##":"Den här staden är fantastisk."
"##actor_good_life##":"Den här staden är inte så illa."
"##lionTamer_need_workers##":"Den här staden behöver mer arbetskraft. Jag undrar om jag kan träna Leo att arbeta mer?"
"##scholar_average_life##":"Den här staden verkar bra."
"##much_plebs##":"Den höga koncentrationen av boende i slumområden i din stad gör att den ser fattig ut."
"##imperial_request_cance_badly_affected##":"Den kejserliga begäran som du nyligen upphävde har skadat din ställning i Rom."
"##high_salary_angers_senate##":"Den löjligt höga lön du betalar till dig själv upprör senaten. Hela Rom talar om din öppna girighet."
"##more_salary_dispeasure_senate##":"Den lön som du betalar dig själv, och som vida överskrider din rang, är en källa till missnöje i Rom."
"##new_governor##":"Den nya guvernören"
"##market_kid_say_1##":"Den tjocka damen bad mig bära detta och följa efter henne."
"##bad_house_quality##":"Den totala kvaliteten på byggnaderna i din stad inverkar negativt på denna ställning."
"##people##":"denarer"
"##peoples##":"denarer"
"##person##":"denarer"
"##dn_collected_this_year##":"denarer har betalats hittills i år"
"##dn_per_month##":"denarer per månad"
"##5_entertainment_access##":"Denna boning har begränsad tillgång till underhållning"
"##6_entertainment_access##":"Denna boning har god tillgång till underhållning"
"##1_entertainment_access##":"Denna boning har knappt tillgång till underhållning"
"##3_entertainment_access##":"Denna boning har mycket begränsad tillgång till underhållning"
"##7_entertainment_access##":"Denna boning har mycket god tillgång till underhållning"
"##4_entertainment_access##":"Denna boning har rimlig tillgång till underhållning"
"##9_entertainment_access##":"Denna boning har tillgång till all underhållning som kan önskas"
"##awesome_entertainment_access##":"Denna boning har tillgång till flera platser för underhållning"
"##8_entertainment_access##":"Denna boning har utmärkt tillgång till underhållning"
"##2_entertainment_access##":"Denna boning har viss tillgång till underhållning"
"##house_evolves_at##":"Denna boning kommer snart att utvecklas och få bättre status, som ett resultat av de förbättrade lokala villkoren."
"##no_space_for_evolve##":"Denna boning skulle kunna få ännu högre status om den hade mer utrymme att expandera."
"##lumber_mill_need_some_workers##":"Denna brädgård arbetar inte med maximal kapacitet. Som resultat kommer timmerproduktionen att bli något långsammare."
"##lumber_mill_full_work##":"Denna brädgård har alla anställda den behöver. Den arbetar fullt ut med att såga timmer."
"##lumber_mill_no_workers##":"Denna brädgård har inga anställda. Produktionen har upphört."
"##bridge_extends_city_area##":"Denna bro ger oss mer mark, men ger fri passage både för medborgare och fiender!"
"##well_haveno_houses_inarea##":"Denna brunn är överflödig för tillfället, eftersom det inte finns några hus inom dess serviceområde."
"##trouble_most_fire##":"Denna byggnad är en brandfara"
"##trouble_no_damage##":"Denna byggnad är i perfekt strukturellt skick"
"##trouble_too_far_from_water##":"Denna byggnad är inte intill vatten!"
"##very_high_damage_risk##":"Denna byggnad är ostadig, och kommer sannolikt att falla samman snart"
"##trouble_some_fire##":"Denna byggnad har brandrisk"
"##middle_file_risk##":"Denna byggnad har en viss brandrisk"
"##working_have_bad_labor_access##":"Denna byggnad har för närvarande dålig tillgång till arbetskraft"
"##working_have_good_labor_access##":"Denna byggnad har för närvarande god tillgång till arbetskraft"
"##working_have_no_labor_access##":"Denna byggnad har för närvarande ingen tillgång till arbetskraft"
"##working_have_very_little_labor_access##":"Denna byggnad har för närvarande mycket liten tillgång till arbetskraft"
"##working_have_awesome_labor_access##":"Denna byggnad har för närvarande utmärkt tillgång till arbetskraft"
"##working_have_some_labor_access##":"Denna byggnad har för närvarande viss tillgång till arbetskraft"
"##trouble_low_fire_risk##":"Denna byggnad har ingen brandrisk"
"##trouble_most_damage##":"Denna byggnad har många strukturella brister och sprickor"
"##very_low_damage_risk##":"Denna byggnad har vissa strukturella brister"
"##moment_fire_risk##":"Denna byggnad kan fatta eld när som helst!"
"##trouble_need_road_access##":"Denna byggnad kräver åtkomst till väg"
"##need_grape##":"Denna byggnad kräver druvor"
"##need_iron_for_work##":"Denna byggnad kräver järnmalm"
"##need_clay_pit##":"Denna byggnad kräver lera"
"##trouble_need_olive##":"Denna byggnad kräver oliver"
"##trouble_need_timber##":"Denna byggnad kräver timmer"
"##trouble_have_damage##":"Denna byggnad löper en liten risk att kollapsa"
"##trouble_some_damage##":"Denna byggnad löper försumbar risk att kollapsa"
"##some_low_fire_risk##":"Denna byggnad utgör en försumbar brandrisk"
"##meat_farm_need_some_workers##":"Denna farm är underbemannad. Svinen har små kullar, som växer långsamt."
"##meat_farm_patrly_workers##":"Denna farm arbetar inte med maximal kapacitet. Som resultat kommer köttproduktionen att bli något mindre."
"##meat_farm_full_work##":"Denna farm har alla anställda den behöver, och dess djurstam är fet och stor."
"##meat_farm_no_workers##":"Denna farm har inga anställda, och alla djuren har flytt eller dött."
"##need_reservoir_for_work##":"Denna fontän fungerar inte eftersom den inte ligger i ett område som täcks av rörledningar från en fungerande reservoar."
"##fountain_not_work##":"Denna fontän fungerar inte eftersom det inte finns tillräckligt med arbetare för att driva den."
"##fountain_will_soon_be_hooked##":"Denna fontän väntar på att anslutas till det underjordiska rörledningsnätet."
"##fig_farm_need_some_workers##":"Denna fruktträdgård är underbemannad. Den producerar mindre frukt än vad den borde."
"##fig_farm_full_work##":"Denna fruktträdgård har alla anställda den behöver. Träden dignar av mogen frukt."
"##fig_farm_no_workers##":"Denna fruktträdgård har inga anställda. Produktionen har upphört."
"##fig_farm_patrly_workers##":"Denna fruktträdgård utnyttjar inte maximal kapacitet. Som resultat kommer fruktproduktionen att gå långsammare."
"##reservoir_info##":"Denna gigantiska cistern innehåller rent dricksvatten, som distribueras via rör av lera över en stor radie i staden. Akvedukter kan länka samman reservoarerna över stora avstånd."
"##trouble_hippodrome_full_work##":"Denna hippodrom har ofta spännande kapplöpningar, som ger mycket nöje åt lokalbefolkningen."
"##trouble_hippodrome_no_charioters##":"Denna hippodrom kör inga kapplöpningar. Den behöver körsvenner."
"##inland_lake_text##":"Denna insjö saknar kontakt med havet"
"##clinic_no_workers##":"Denna klinik används inte, och är därför värdelös för lokalsamhället."
"##clinic_full_work##":"Denna klinik används, och betjänar lokalsamhället."
"##wheat_farm_need_some_workers##":"Denna lantgård är underbemannad. Arbetarna kan inte så alla de fält som finns."
"##vegetable_farm_need_some_workers##":"Denna lantgård är underbemannad. Vissa av dess grönsaker kommer att ruttna på åkern."
"##wheat_farm_patrly_workers##":"Denna lantgård arbetar under sin maximala kapacitet. Fler arbetare skulle öka produktiviteten."
"##wheat_farm_full_work##":"Denna lantgård har alla anställda det behöver. Den får maximum avkastning på sin areal."
"##vegetable_farm_full_work##":"Denna lantgård har alla anställda det behöver. Grönsaker växer här i överflöd."
"##olive_farm_no_workers##":"Denna lantgård har inga anställda. Inget har planterats."
"##vegetable_farm_no_workers##":"Denna lund har inga anställda. Produktionen har upphört."
"##wheat_farm_no_workers##":"Denna lantgård har inga anställda. Jorden ligger i träda."
"##vegetable_farm_patrly_workers##":"Denna lantgård utnyttjar inte maximal kapacitet. Därför kommer grönsaksproduktionen att gå något långsammare."
"##legion_haveho_soldiers_and_barracks##":"Denna legion har för närvarande inga soldater. Den existerar bara till namnet och utan förläggningar i staden kan den inte ta emot några nya trupper."
"##legion_haveho_soldiers##":"Denna legion har för närvarande inga soldater. Den existerar bara till namnet. Endast när nyligen utbildade trupper anländer från förläggningarna kommer den att förvandlas till en stridande enhet."
"##olive_farm_patrly_workers##":"Denna lund är underbemannad. Det tar längre tid att plocka oliverna än vad det borde."
"##olive_farm_full_work##":"Denna lund har alla anställda den behöver. Trädgrenarna dignar med tunga lass av oliver."
"##olive_farm_need_some_workers##":"Denna lund utnyttjar inte maximal kapacitet. Olivproduktionen kan bli bättre med fler arbetare."
"##market_full_work##":"Denna marknad används"
"##market_no_workers##":"Denna marknad används inte, och levererar inga produkter till lokalsamhället."
"##market_search_food_source##":"Denna marknad har köpmän men de söker för närvarande efter en källa till livsmedel som kan säljas."
"##vinard_need_some_workers##":"Denna odling är underbemannad. Det tar längre tid att producera druvor än vad det borde."
"##vinard_full_work##":"Denna odling har alla anställda den behöver. Vinrankorna är tunga med stora, saftiga druvor."
"##vinard_no_workers##":"Denna odling har inga anställda. Produktionen har upphört."
"##vinard_patrly_workers##":"Denna odling utnyttjar inte maximal kapacitet. Som resultat kommer druvproduktionen att bli mindre."
"##oil_workshop_full_work##":"Denna olivpress är fullt bemannad och producerar rikliga mängder olja av hög kvalitet."
"##oil_workshop_patrly_workers##":"Denna olivpress är underbemannad och producerar oljan mycket långsammare än vad den borde."
"##oil_workshop_need_some_workers##":"Denna olivpress behöver fler arbetare för att nå sin fulla potential för oljeproduktion."
"##oil_workshop_no_workers##":"Denna olivpress har inga anställda och kommer inte att producera olja."
"##oil_workshop_need_resource##":"Denna olivpress kommer inte att producera olja utan leverans av oliver, från ett magasin eller från en lantgård."
"##mopup_formation_text##":"Denna ordning är det effektivaste sättet att hantera resterna av en besegrad armé."
"##province_has_peace_a_short_time##":"Denna provins har haft fred en kort tid, men dina invånare känner sig fortfarande inte helt säkra. Fler fredsår kommer att förbättra detta."
"##this_province_feels_peaceful##":"Denna provins känns förhållandevis säker, en känsla som kan förbättras med tiden."
"##reservoir_no_water##":"Denna reservoar fungerar inte eftersom den inte ligger intill vatten eller inte är ansluten till en annan reservoar via akvedukter."
"##school_no_workers##":"Denna skola används inte, och är värdelös för lokalsamhället."
"##school_full_work##":"Denna skola används, och barnen i stadsdelen är läskunniga och vältaliga."
"##weapons_workshop_need_some_workers##":"Denna smedja är underbemannad, och det tar längre tid att producera vapen än vad det borde."
"##weapons_workshop_full_work##":"Denna smedja har alla anställda den behöver, den arbetar fullt ut med att producera vapen."
"##weapons_workshop_patrly_workers##":"Denna smedja utnyttjas inte till maximal kapacitet. Vapenproduktionen kommer att gå något långsammare än vad den borde."
"##marketBuyer_average_life##":"Denna stad är egentligen inte så illa."
"##priest_average_life##":"Denna stad är en hygglig plats att bo på."
"##prefect_need_workers##":"Denna stad är i desperat behov av arbetare!"
"##priest_low_entertainment##":"Denna stad är så tråkig. Även en präst tycker om gladiatorspel då och då."
"##theater_no_have_any_shows##":"Denna teater har sällan några uppsättningar. Den behöver riktiga skådespelare för att kunna erbjuda underhållning."
"##theater_full_work##":"Denna teater sätter för närvarande upp pjäser med lokala aktörer, som vanligen drar stor publik."
"##garden_info##":"Denna trevliga plats skänker medborgarna avkoppling från stadens buller, värme och smuts genom en sval oas av grönska. Alla vill ha en trädgård intill sitt hus."
"##weapons_workshop_no_workers##":"Denna vapenfabrik har inga anställda. Produktionen har upphört."
"##furniture_workshop_no_workers##":"Denna verkstad har inga anställda. Produktionen har upphört."
"##weapons_workshop_need_resource##":"Denna verkstad kräver leverans av järn, från ett magasin eller från ett malmbrott, för att producera vapen."
"##wine_workshops_need_some_workers##":"Denna vingård är underbemannad och det tar mycket längre tid att producera vin än vad det borde."
"##wine_workshop_full_work##":"Denna vingård har alla anställda den behöver och arbetar fullt ut med att producera vin."
"##wine_workshop_no_workers##":"Denna vingård har inga anställda. Produktionen har upphört."
"##wine_workshop_need_resource##":"Denna vingård kan inte producera vin förrän den får en leverans av druvor från ett magasin eller en druvodling."
"##wine_workshops_patrly_workers##":"Denna vingård utnyttjar inte full kapacitet. Vinproduktionen något långsammare än vad den borde vara."
"##enemies_hard_to_me##":"Denne soldat är för stark för mig!"
"##engineer_have_trouble_buildings##":"Dessa byggnader är i dåligt skick. Jag kom precis i rätt tid."
"##this_fire_can_spread##":"Dessa eldsvådor sprider sig om du inte snabbt hejdar dem."
"##taxCollector_very_little_tax##":"Dessa hus betalar så lite skatt att det är slöseri med tiden."
"##these_rift_info##":"Dessa klyftor har orsakats av jordbävningar. De kan inte passeras eller fyllas."
"##marketBuyer_return##":"Dessa korgar är så tunga! Jag har med mig färska varor till min marknad."
"##collapsed_ruins_info##":"Dessa spillror av gamla byggnader gör marken mindre åtråvärd."
"##these_goods_import_only##":"Dessa varor finns endast tillgängliga via import"
"##balance_between_migration##":"Det är lika många som kommer till, respektive lämnar staden"
"##lion_pit_work##":"Det är med nöje vi tillkännager att vi, med full sysselsättning, kan leverera upp till fyra nya lejon varje månad."
"##gladiator_pit_full_work##":"Det är med nöje vi tillkännager att vi, med full sysselsättning, utbildar upp till fyra nya gladiatorer varje månad."
"##lionTamer_high_workless##":"Det är stor arbetslöshet här."
"##massilia_preview_mission##":"Det enda vattnet finns i oasen. Detsamma gäller tyvärr för odlingsbar mark. Reservoarer och lantgårdar konkurrerar om samma utrymme. Använd det med förstånd."
"##emperor_send_money_to_you_nearest_time##":"Det faktum att kejsaren nyligen måste ingripa för att rädda dig skadar allvarligt din stads rykte om välstånd."
"##amazing_prosperity_this_city##":"Det fantastiska välståndet i den här staden är det stora samtalsämnet i Rom!"
"##shipyard_notneed_ours_boat##":"Det finns för närvarande inga fiskehamnar som behöver våra båtar."
"##actor_need_workers##":"Det finns helt enkelt inte tillräckligt med arbetare i staden."
"##need_trainee_charioteer##":"Det finns inga kapplöpningsvagnar i din hippodrom. Anskaffning av sådana skulle avsevärt förbättra villkoren för befolkningen, som ivrigt söker mer underhållning."
"##prefect_so_hungry##":"Det finns inte nog med mat i staden. Det ökar brottsligheten."
"##marketBuyer_so_hungry##":"Det finns inte tillräckligt med livsmedel här. Hur ska jag kunna försörja mig?"
"##vegetable_farm_bad_work##":"Det finns knappt några anställda för att underhålla jordbruket, de få grönsakerna kommer att bli offer för insekter."
"##meat_farm_bad_work##":"Det finns knappt några anställda vid den här farmen, djurantalet e lågt och växer extremt långsamt."
"##advchief_low_crime##":"Det finns lite brottslighet här, ingenting allvarligt."
"##wheat_farm_bad_work##":"Det finns mycket få jordbruksarbetare här. Som resultat är veteproduktionen långsam."
"##olive_farm_slow_work##":"Det finns mycket få människor som arbetar här. Som resultat är olivproduktionen långsam."
"##vinard_bad_work##":"Det finns nästan inga anställda på denna vinodling. Som resultat kommer mycket få druvor att klara sig till skörden."
"##lumber_mill_bad_work##":"Det finns nästan inga skogsarbetare, produktionen står nästan helt still."
"##scholar_need_workers##":"Det finns så få arbetare att någon till och med erbjöd mig jobb."
"##cartSupplier_average_life##":"Det här är en bra stad. Folk tycker om att bo här."
"##small_colloseum_show##":"Det krävs fler spektakel i dina colosseum! Genom att förse dem med gladiatorer eller lejon förbättras underhållningen i delar av staden."
"##barber_need_workers##":"Det saknas många arbetare här."
"##engineering_post_need_some_workers##":"Det tar en eller två dagar innan våra utarbetade ingenjörer är tillbaka på gatorna."
"##road_to_distant_region##":"Detta är den väg som leder till rikets utposter. Det är en kejserlig huvudväg, som måste hållas öppen längs hela sin sträckning."
"##doctor_average_life##":"Detta är en fantastisk stad."
"##peaceful_crime_risk##":"Detta är en fridfull stadsdel."
"##marketBuyer_gods_angry##":"Detta är en hednisk plats. Ståthållaren har ingen respekt för gudarna."
"##this_lawab_province_become_very_peacefull##":"Detta är en laglydig provins som med tiden kan bli mycket fredlig."
"##cartSupplier_good_life##":"Detta är en magnifik stad."
"##very_low_crime_risk##":"Detta är en mycket laglydig stadsdel, ingen brottslighet alls"
"##prefect_good_life##":"Detta är en underbar plats att bo på."
"##averange_crime_risk##":"Detta är ett område med hög brottslighet. De boende är missnöjda, och gatorna är farliga"
"##few_crime_risk##":"Detta är ett område med låg brottslighet, men vissa boende har klagat"
"##overall_city_become_a_sleepy_province##":"Detta är på det hela taget en provins med få verkliga hot - precis så som invånarna vill ha det!"
"##this_is_ruins##":"Detta är spillrorna från byggnaden som nämns ovan. Förfallna platser gör inte att området ser vackrare ut."
"##road_from_rome##":"Detta är vägen till Rom. Immigranterna anländer från denna punkt. Därför är det viktigt att vägen hålls öppen. Även köpmän passerar genom din provins längs denna kejserliga huvudväg."
"##library_full_work##":"Detta bibliotek används. Dess hyllor är fyllda med skriftrullar med lärdom."
"##iron_mine_patrly_workers##":"Detta brott är underbemannat. Det tar längre tid än normalt att producera järnet."
"##quarry_full_work##":"Detta brott har alla anställda det behöver, det arbetar fullt ut med att producera marmor."
"##iron_mine_full_work##":"Detta brott har alla anställda det behöver, och arbetar fullt ut med att producera järn."
"##quarry_no_workers##":"Detta brott har inga anställda. Produktionen har upphört."
"##iron_mine_no_workers##":"Detta brott har inga anställda. Produktionen har upphört."
"##iron_mine_need_some_workers##":"Detta brott utnyttjar inte maximal kapacitet. Malmbrytningen skulle vara mycket effektivare med fler arbetare."
"##quarry_need_some_workers##":"Detta brott utnyttjar inte maximal kapacitet. Som resultat kommer marmorproduktionen att bli något mindre."
"##colloseum_no_workers##":"Detta colosseum är stängt. Utan anställda är det värdelöst som rekreationsanläggning."
"##trouble_colloseum_full_work##":"Detta colosseum har både gladiatorkamp och lejonkamper, till lokalsamhällets stora nöje."
"##trouble_colloseum_have_only_lions##":"Detta colosseum har djurkamp, med lejon från lokala handelsmän. Den skulle också kunna anlita gladiatorer för kamp man mot man."
"##trouble_colloseum_have_only_gladiatros##":"Detta colosseum har gladiatorkamp för lokalbefolkningen. Lejon skulle ge mer variation till dödskamperna."
"##trouble_colloseum_no_shows##":"Detta colosseum har inga föreställningar. Det behövs gladiatorer och lejon för att locka publik."
"##fort_has_been_cursed_by_mars##":"Detta fort har förbannats av Mars. Det kommer att dröja innan några soldater vågar sig tillbaka hit."
"##house_not_registered_for_taxes##":"Detta hus befinner sig i en region utan skatteadministration, och betalar därför ingen skatt"
"##religion_access_1_temple##":"Detta hus har endast tillgång till ett tempel för en enda gud"
"##education_have_no_access##":"Detta hus har ingen grundläggande tillgång till skolor eller bibliotek"
"##colosseum_no_access##":"Detta hus har ingen tillgång till ett colosseum"
"##house_have_not_food##":"Detta hus har inget livsmedelsförråd"
"##house_no_troubles_with_food##":"Detta hus har inget problem med att skaffa den mat som krävs för att överleva"
"##warning_amphitheater_access##":"Detta hus har inte passerats av en gladiator på ett tag. Det kommer snart att förlora tillgång till amfiteater"
"##warning_hippodrome_access##":"Detta hus har inte passerats av en körsven på ett tag. Det kommer snart att förlora tillgång till hippodrom"
"##warning_colloseum_access##":"Detta hus har inte passerats av en lejontämjare på ett tag. Det kommer snart att förlora tillgång till colosseum"
"##warning_theater_access##":"Detta hus har inte passerats av en skådespelare på ett tag. Det kommer snart att förlora tillgången till teater"
"##library_no_access##":"Detta hus har inte tillgång till bibliotek"
"##no_academy_access##":"Detta hus har inte tillgång till en högskola"
"##doctor_no_access##":"Detta hus har inte tillgång till en klinik"
"##theater_no_access##":"Detta hus har inte tillgång till en teater"
"##hospital_no_access##":"Detta hus har inte tillgång till ett sjukhus"
"##hippodrome_no_access##":"Detta hus har inte tillgång till hippodromen"
"##school_no_access##":"Detta hus har inte tillgång till någon skola"
"##religion_no_access##":"Detta hus har inte tillgång till några tempel eller orakel"
"##house_food_only_for_month##":"Detta hus har matförråd som åtminstone kommer att räcka under den kommande månaden"
"##awesome_amphitheater_access##":"Detta hus har tillgång till amfiteater"
"##library_full_access##":"Detta hus har tillgång till bibliotek"
"##awesome_colloseum_access##":"Detta hus har tillgång till colosseum"
"##awesome_doctor_access##":"Detta hus har tillgång till en klinik"
"##religion_access_full##":"Detta hus har tillgång till ett orakel, och till tempel för alla gudar"
"##hippodrome_full_access##":"Detta hus har tillgång till hippodrom"
"##education_have_academy_access##":"Detta hus har tillgång till högskola"
"##hospital_full_access##":"Detta hus har tillgång till sjukhus"
"##school_full_access##":"Detta hus har tillgång till skola"
"##education_have_school_or_library_access##":"Detta hus har tillgång till skola eller bibliotek"
"##education_have_school_library_access##":"Detta hus har tillgång till skola och bibliotek"
"##education_full_access##":"Detta hus har tillgång till skola, bibliotek och högskola"
"##theater_full_access##":"Detta hus har tillgång till teater"
"##religion_access_2_temple##":"Detta hus har tillgång till tempel för 2 olika gudar"
"##religion_access_3_temple##":"Detta hus har tillgång till tempel för 3 olika gudar"
"##religion_access_4_temple##":"Detta hus har tillgång till tempel för 4 olika gudar"
"##religion_access_5_temple##":"Detta hus har tillgång till tempel för alla gudarna"
"##missing_college##":"Detta hus kan inte utvecklas, eftersom dess redan utmärkta tillgång till utbildning måste förbättras genom tillgång till en högskola."
"##missing_school##":"Detta hus kan inte utvecklas, eftersom dess tillgång till utbildning måste förbättras genom tillgång till en skola."
"##missing_library##":"Detta hus kan inte utvecklas, eftersom dess tillgång till utbildning måste förbättras genom tillgång till ett bibliotek."
"##missing_second_religion##":"Detta hus kan inte utvecklas, eftersom det endast har tillgång till tempel för en enda gud. I takt med att dess invånare kommer upp sig i världen kommer de att vilja ägna mer tid åt att tillbe andra gudar."
"##missing_third_religion##":"Detta hus kan inte utvecklas, eftersom det endast har tillgång till tempel för två gudar. I takt med att dess invånare kommer upp sig i världen kommer de att vilja ägna mer tid åt att tillbe andra gudar."
"##missing_doctor_or_hospital##":"Detta hus kan inte utvecklas, eftersom det i stort sett saknar tillgång till sjukvård. Det saknar tillgång till både klinik och sjukhus."
"##missing_entertainment##":"Detta hus kan inte utvecklas, eftersom det inte finns någon underhållning i området."
"##missing_entertainment_also##":"Detta hus kan inte utvecklas, eftersom det inte finns tillräckligt med underhållning i området."
"##missing_barber##":"Detta hus kan inte utvecklas, eftersom det inte har någon lokal tillgång till en barberare."
"##missing_market##":"Detta hus kan inte utvecklas, eftersom det inte har tillgång till en lokal marknad."
"##missing_water##":"Detta hus kan inte utvecklas, eftersom det inte har tillgång till ens den mest primitiva vattenförsörjning."
"##missing_bath##":"Detta hus kan inte utvecklas, eftersom det inte har tillgång till ett lokalt badhus."
"##missing_school_or_library##":"Detta hus kan inte utvecklas, eftersom det inte har tillgång till grundläggande utbildningsmöjligheter vare sig från skola eller bibliotek."
"##missing_religion##":"Detta hus kan inte utvecklas, eftersom det inte har tillgång till några lokala möjligheter till religionsutövning."
"##missing_fountain##":"Detta hus kan inte utvecklas, eftersom det inte har tillgång till ren vattentillförsel från en fontän."
"##missing_entertainment_amph##":"Detta hus kan inte utvecklas, eftersom det knappt finns någon underhållning i området."
"##missing_second_food##":"Detta hus kan inte utvecklas, eftersom det krävs en till typ av livsmedel, som levereras från en lokal marknad, för att förmå mer välbärgade att flytta in."
"##missing_third_food##":"Detta hus kan inte utvecklas, eftersom det krävs en tredje typ av livsmedel, som levereras från en lokal marknad, för att förmå patricierklasserna att flytta in."
"##missing_food##":"Detta hus kan inte utvecklas, eftersom det måste ha leveranser av livsmedel från en lokal marknad."
"##missing_doctor##":"Detta hus kan inte utvecklas, eftersom det vill ha bättre möjligheter till sjukvård. Det finns lokal tillgång till ett sjukhus men det behövs en klinik i närheten."
"##missing_hospital##":"Detta hus kan inte utvecklas, eftersom det vill ha bättre möjligheter till sjukvård. Klinikernas täckning är bra men det saknas lokal tillgång till ett sjukhus."
"##missing_entertainment_need_more##":"Detta hus kan inte utvecklas, eftersom det visserligen finns god underhållning i området, men inte tillräckligt varierat utbud."
"##missing_entertainment_patrician##":"Detta hus kan inte utvecklas, eftersom det visserligen finns utmärkt underhållning i området, men det är trångt och utbudet är inte tillräckligt varierat för de kräsna patricierna."
"##missing_entertainment_colloseum##":"Detta hus kan inte utvecklas, eftersom det visserligen finns viss underhållning i området, men inte tillräckligt."
"##missing_pottery##":"Detta hus kan inte utvecklas. Det behöver leveranser av krukor från sin lokala marknad innan förmögnare medborgarklasser kommer att flytta in."
"##missing_oil##":"Detta hus kan inte utvecklas. Det behöver oljeleveranser från sin lokala marknad innan mer välmående medborgarklasser kommer att flytta in."
"##missing_furniture##":"Detta hus kan inte utvecklas. Det behöver tillgång till möbelleveranser från sin lokala marknad innan mer välmående medborgarklasser kommer att flytta in."
"##missing_wine##":"Detta hus kan inte utvecklas. Det behöver tillgång till vinleveranser från sin lokala marknad innan mer välmående medborgarklasser kommer att flytta in."
"##missing_food_from_market##":"Detta hus kan inte utvecklas. Det har visserligen tillgång till en lokal marknad, men marknaden själv har svårt att få livsmedelsleveranser."
"##missing_second_wine##":"Detta hus kan inte utvecklas. Det krävs en vinsort till för att tillfredsställa de sysslolösa patriciernas dekadenta livsstil. Öppna en ny handelsväg, eller tillverka ditt eget vin."
"##house_have_some_food##":"Detta hus kommer snart att äta upp sitt begränsade livsmedelsförråd"
"##missing_doctor__degrade##":"Detta hus kommer snart att förfalla, eftersom dess möjligheter till hälsovård skurits ned. Det finns lokal tillgång till ett sjukhus men det är svårt att hitta en klinik."
"##missing_hospital_degrade##":"Detta hus kommer snart att förfalla, eftersom dess tillgång till hälsovård har skurits ned. Tillgången till kliniker är god men det finns inga lokala sjukhus."
"##missing_third_food_degrade##":"Detta hus kommer snart att förfalla, eftersom det endast har tillgång till 2 typer av livsmedel från sin lokala marknad. Detta avskräcker patricierklasserna."
"##missing_second_food_degrade##":"Detta hus kommer snart att förfalla, eftersom det endast har tillgång till en enda typ av livsmedel från sin lokala marknad. Detta avskräcker de välbärgade klasserna."
"##missing_religion_degrade##":"Detta hus kommer snart att förfalla, eftersom det har förlorat all tillgång till lokala religiösa byggnader."
"##missing_school_or_library_degrade##":"Detta hus kommer snart att förfalla, eftersom det har förlorat alla grundläggande utbildningsmöjligheter från en skola eller ett bibliotek."
"##missing_barber_degrade##":"Detta hus kommer snart att förfalla, eftersom det har förlorat tillgången till barberare."
"##missing_bath_degrade##":"Detta hus kommer snart att förfalla, eftersom det har förlorat tillgången till sitt badhus."
"##missing_furniture_degrade##":"Detta hus kommer snart att förfalla, eftersom det har slut på möbler och dess lokala marknad har ett sporadiskt utbud."
"##missing_oil_degrade##":"Detta hus kommer snart att förfalla, eftersom det har slut på oljan och dess lokala marknad har ett sporadiskt utbud."
"##missing_wine_degrade##":"Detta hus kommer snart att förfalla, eftersom det har slut på vin och dess lokala marknad har ett sporadiskt utbud."
"##missing_entertainment_degrade##":"Detta hus kommer snart att förfalla, eftersom det knappast finns någon underhållning i området."
"##missing_food_degrade##":"Detta hus kommer snart att förfalla. Det har visserligen tillgång till en marknad, men marknaden själv har svårt att få livsmedelsleveranser."
"##missing_fountain_degrade##":"Detta hus kommer snart att förfalla, eftersom det inte har tillgång till rent vatten från en fontän."
"##missing_doctor_or_hospital_degrade##":"Detta hus kommer snart att förfalla, eftersom det nu har tvivelaktig hälsovård. Det saknas inte bara tillgång till en klinik, utan även tillgången till sjukhus är dålig."
"##missing_water_degrade##":"Detta hus kommer snart att förfalla, eftersom det saknar tillgång till även den enklaste vattenförsörjning."
"##low_desirability_degrade##":"Detta hus kommer snart att förfalla. Den sjunkande efterfrågan på boende i detta område drar ner det."
"##missing_third_religion_degrade##":"Detta hus kommer snart att förfalla. Dess tidigare utmärkta religiösa möjligheter har reducerats, och det har nu endast tillgång till tempel för två gudar."
"##missing_college_degrade##":"Detta hus kommer snart att förfalla. Dess tidigare utmärkta tillgång till utbildning har försämrats, eftersom det har förlorat tillgången till sin högskola."
"##missing_second_religion_degrade##":"Detta hus kommer snart att förfalla. Dess tillgång till lokala religiösa byggnader har reducerats till endast ett tempel för en enda gud."
"##missing_school_degrade##":"Detta hus kommer snart att förfalla. Dess tillgång till utbildning har försämrats, eftersom det har förlorat tillgång till sin skola."
"##missing_library_degrade##":"Detta hus kommer snart att förfalla. Dess tillgång till utbildning har försämrats, eftersom det har förlorat tillgång till sitt bibliotek."
"##missing_entertainment_also_degrade##":"Detta hus kommer snart att förfalla. Det finns god underhållning i området, men inte tillräckligt varierat utbud."
"##missing_entertainment_colloseum_degrade##":"Detta hus kommer snart att förfalla. Det finns utmärkt underhållning i området, men det är trångt och utbudet är inte tillräckligt varierat för de kräsna patricierna."
"##missing_entertainment_amph_degrade##":"Detta hus kommer snart att förfalla. Det finns viss underhållning i området, men inte tillräckligt."
"##missing_market_degrade##":"Detta hus kommer snart att förfalla. Det har förlorat tillgången till en marknad."
"##missing_pottery_degrade##":"Detta hus kommer snart att förfalla. Det har inte längre tillgång till krukor, och leveranserna till dess lokala marknad är minst sagt opålitliga."
"##pottery_workshop_need_som_workers##":"Detta krukmakeri är underbemannat och produktionen tar längre tid än normalt."
"##pottery_workshop_need_resource##":"Detta krukmakeri behöver leveranser av lera, från ett magasin eller från ett lertag, för att kunna producera krukor."
"##pottery_workshop_full_work##":"Detta krukmakeri har alla anställda det behöver. Det arbetar fullt ut med att producera krukor."
"##pottery_workshop_patrly_workers##":"Detta krukmakeri utnyttjar inte maximal kapacitet. Som resultat kommer krukproduktionen att gå långsammare."
"##desirability_pretty_area##":"Detta land är ett eftertraktat område, vad gäller dina medborgare"
"##clear_land_text##":"Detta landområde kan byggas på efter behov. Det ger fri passage både åt egna soldater och åt fiendesoldater."
"##triumphal_arch_info##":"Detta magnifika byggnadsverk är tillägnat Roms historiska segrar över sina fiender. Inget kan ge högre status."
"##dangerous_crime_risk##":"Detta område är farligt."
"##water_srvc_well##":"Detta område har tillgång till dricksvatten"
"##water_srvc_fountain_and_well##":"Detta område har tillgång till en reservoar via rörledning och dricksvatten från en brunn eller fontän"
"##water_srvc_reservoir##":"Detta område har tillgång till en reservoar via rörledning, vilket gör att fontäner och badhus fungerar"
"##high_crime_risk##":"Hela detta område är som en jäsande krutdurk! Brottsligheten är epidemisk, och uppror sannolika"
"##hospital_no_workers##":"Detta sjukhus används inte, och är därför värdelöst för lokalsamhället."
"##hospital_full_work##":"Detta sjukhus används, och betjänar lokalsamhället."
"##furniture_workshop_need_some_workers##":"Detta snickeri är underbemannat, och det tar längre tid att producera möbler än vad det borde."
"##furniture_workshop_need_resource##":"Detta snickeri behöver leverans av virke från ett magasin eller från en brädgård för att kunna producera möbler."
"##furniture_workshop_full_work##":"Detta snickeri har full sysselsättning, och arbetar fullt ut med att producera möbler."
"##furniture_workshop_patrly_workers##":"Detta snickeri har lediga platser. Möbelproduktionen blir effektivare när de fyllts."
"##big_fest_description##":"Din 2 dagars festival för din valda gud är slut. Ditt folk respekterar dig."
"##lugdunum_win_text##":"Din behandling av gallerna i Lugdunum och den sköna stadens prakt bådar väl för Roms expansion i den norra vildmarken. Bra gjort!"
"##capua_win_text##":"Din förmåga att styra imponerar på mig. Många ståthållares karriärer gäckas när jag ber dem bygga den första kolonin. Ledare som du garanterar Rom en framtid. Kan du upprepa dina framgångar eller var det bara tur?"
"##broke_empiretax_with2years_warning##":"Din fortsatta oförmåga att lämna tribut till Rom skadar ditt rykte."
"##trade_advisor_blocked_timber_production##":"Din handelsrådgivare har stoppat all avverkning."
"##trade_advisor_blocked_grape_production##":"Din handelsrådgivare har stoppat all druvodling."
"##trade_advisor_blocked_fruit_production##":"Din handelsrådgivare har stoppat all fruktodling."
"##trade_advisor_blocked_vegetable_production##":"Din handelsrådgivare har stoppat all grönsaksodling."
"##trade_advisor_blocked_meat_production##":"Din handelsrådgivare har stoppat all köttproduktion."
"##trade_advisor_blocked_pottery_production##":"Din handelsrådgivare har stoppat all kruktillverkning."
"##trade_advisor_blocked_iron_production##":"Din handelsrådgivare har stoppat all malmbrytning."
"##trade_advisor_blocked_marble_production##":"Din handelsrådgivare har stoppat all marmorbrytning."
"##trade_advisor_blocked_furniture_production##":"Din handelsrådgivare har stoppat all möbeltillverkning."
"##trade_advisor_blocked_olive_production##":"Din handelsrådgivare har stoppat all olivodling."
"##trade_advisor_blocked_oil_production##":"Din handelsrådgivare har stoppat all oljeproduktion."
"##trade_advisor_blocked_weapon_production##":"Din handelsrådgivare har stoppat all vapenproduktion."
"##trade_advisor_blocked_wheat_production##":"Din handelsrådgivare har stoppat all veteodling."
"##trade_advisor_blocked_wine_production##":"Din handelsrådgivare har stoppat all vinproduktion."
"##trade_advisor_blocked_clay_production##":"Din handelsrådgivare har stoppat alla lertag."
"##not_enought_place_for_legion##":"Din legion har de fort som krävs"
"##playerarmy_gone_to_location##":"Din legion marscherar för att befria en stad från riket"
"##playerarmy_gone_to_home##":"Din legion på återtåg till din stad"
"##healthadv_noproblem_small_city##":"Din lilla bosättning har ännu inga hälsoproblem att rapportera."
"##request_failed##":"Din nyligen visade oförmåga eller ovilja att utföra en kejserlig begäran har skadat din ställning i Rom en aning."
"##broke_empiretax_warning##":"Din oförmåga att betala tribut till Rom utmålar din stad som misslyckad."
"##your_favor_is_dropping_catch_it##":"Din popularitet i Rom minskar. Du måste fånga Caesars intresse på ett eller annat sätt!"
"##your_province_quiet_and_secure##":"Din provins lugna och säkra tillvaro har blivit legendarisk. Andra ståthållare planerar förmodligen att dra sig tillbaka hit!"
"##cant_calc_prosperity##":"Din stad är ny. Vi har inte haft möjlighet att bedöma ditt välstånd än!"
"##city_has_runout_money##":"Din stad har inga pengar kvar. Caesar har gått med på att ge dig mer, men han kommer inte vara så generös nästa gång. Exportera varor för att generera mer inkomst till din stad."
"##1000_citizens_in_city##":"Din stads population har nått 1.000 invånare för första gången."
"##10000_citizens_in_city##":"Din stads population har nått 10.000 invånare för första gången."
"##100_citizens_in_city##":"Din stads population har nått 100 invånare för första gången."
"##15000_citizens_in_city##":"Din stads population har nått 15.000 invånare för första gången."
"##2000_citizens_in_city##":"Din stads population har nått 2.000 invånare för första gången."
"##20000_citizens_in_city##":"Din stads population har nått 20.000 invånare för första gången."
"##25000_citizens_in_city##":"Din stads population har nått 25.000 invånare för första gången."
"##3000_citizens_in_city##":"Din stads population har nått 3.000 invånare för första gången."
"##5000_citizens_inc_city##":"Din stads population har nått 5.000 invånare för första gången."
"##500_citizens_in_city##":"Din stads population har nått 500 invånare för första gången."
"##your_favour_unchanged_from_last_year##":"Din ställning är oförändrad sedan förra året."
"##your_favour_increased_from_last_year##":"Din ställning i Rom har förbättrats sedan förra året."
"##your_prosperity_raising##":"Din välståndsställning förbättras."
"##we_produce_less_than_eat##":"Dina invånare äter mer mat än de producerar"
"##this_time_you_city_not_need_religion##":"Dina medborgare är ännu så länge upptagna med andra aspekter på stadslivet. I takt med att staden växer kommer de att vilja ha tillgång till ett stort Tempelutbud."
"##need_temples_for_city##":"Dina medborgare har börjat bli intresserade av religion. Frånvaron av en närliggande gudstjänstplats hindrar stadens utveckling."
"##desirability_indiffirent_area##":"Dina medborgare ser varken positivt eller negativt på detta område"
"##gods_unhappy_text##":"Dina medborgarna tror att gudarna kan bli upprörda. Vissa medborgare har visioner av annalkande katastrofer. Bygg nya tempel och börja fester för deras skull, annars riskerar du att drabbas av deras vrede."
"##distribution_center##":"Distributionscentral"
"##more_0_month_from_festival##":"Ditt folk, somliga fortfarande berusade efter festen, välkomnar din generositet."
"##governor_palace_1_info##":"Ditt hem är en av stadens mest attraktiva adresser."
"##more_12_month_from_festival##":"Ditt invånare är mycket missnöjda med tanken på ännu ett år utan en festival."
"##other##":"Diverse"
"##sldr_daring##":"Djärv"
"##denarii_short##":"dn"
"##donation_is##":"Donationen är"
"##send_money##":"Donera dessa pengar till staden från dina personliga besparingar"
"##donations##":"Donerat"
"##vinard##":"Druvodling"
"##vinard_info##":"Druvorna från dessa vinrankor har odlats särskild för vinframställning. Vingårdarna gör fint vin för dina egna patricier, samt för export."
"##tarsus_win_text##":"Du är på god väg att bli min mest uppskattade undersåte. Din mästerliga förståelse av handeln gjorde Tarsus till precis den stad jag hoppats på. De östliga provinserna är mer lojala i dag, tack vare dig."
"##emperor_anger_text##":"Du avsikligt vägrar skicka mig det jag frågat efter? Eller vill du förnedra mig?"
"##oracle_need_2_cart_marble##":"Du behöver 2 ton marmor för att bygga ett orakel"
"##need_marble_for_large_temple##":"Du behöver 2 ton marmor för att bygga ett stort tempel"
"##low_desirability##":"Du behöver göra området mer attraktivt -kanske genom att anlägga några trädgårdar eller torg."
"##city_loathed_you##":"Du föraktas i hela staden"
"##wrath_of_neptune_failed_description##":"Du har åtdragit mitt vrede. Jag ser fram emot när din stad börjar använda båtar, då kommer hämnden."
"##have_less_library_in_city_0##":"Du har för få bibliotek i din stad. Om du bygger fler förbättras din ställning."
"##have_less_academy_in_city_0##":"Du har för få högskolor i din stad. Om du bygger fler förbättras din ställning."
"##have_less_temple_in_city_0##":"Du har för få religiösa byggnader i din stad. Om du bygger fler förbättras din ställning."
"##have_less_school_in_city_0##":"Du har för få skolor i din stad. Om du bygger fler förbättras din ställning."
"##have_less_theater_in_city_0##":"Du har för få teatrar i din stad. Om du bygger fler förbättras din ställning."
"##legionadv_no_legions##":"Du har inga legioner att leda. Du måste först bygga ett fort"
"##have_no_legions##":"Du har inga legioner att sända"
"##no_culture_building_in_city##":"Du har ingen kultur i din stad, ergo (latin för därför!) har du ingen kulturställning."
"##current_year_notpay_tribute_warning##":"Du har inte betalat tribut detta året. Spara lite pengar i din skattkammare så att du kan göra din årliga betalning."
"##nomoney_for_gift_text##":"Du har inte tillräcklig med personliga besparingar för att kunna betala en gåva till kejsaren. Försök att betala dig själv högre lön!"
"##no_goods_for_request##":"Du har inte tillräckligt med varor i dina handelsmagasin"
"##city_has_runout_money_again##":"Du har slösat med Roms tillgångar. Caesar har ilsket gått med på att låna 5.000 denarii for 12 månader. Du behöver generera pengar från skatt och exportering."
"##can_build_only_one_of_building##":"Du kan endast ha en byggnad av denna typ"
"##tutorial2_win_text##":"Du lär dig snabbt! Nu har du tillräckligt med kunskap för att klara ett riktigt uppdrag. Från och med nu kan du välja vilken riktning din karriär ska ta. Välj en fredligare provins om du vill koncentrera dig på att styra eller en farligare provins om du vill tampas med Roms fiender."
"##need_build_on_cleared_area##":"Måste byggas på avröjt land"
"##edil_salary##":"Edillön på"
"##effciency##":"Effektivitet"
"##egift_egyptian_glassware##":"Egyptiska glasvaror"
"##no_visited_by_taxman##":"Ej fått besök av skatteindrivare. Betalar ej skatt"
"##not_available##":"Ej tillgänglig... ännu!"
"##city_fire_title##":"Eldsvåda i din stad"
"##emigrant##":"Emigrant"
"##wt_emigrant##":"Emigrant"
"##distant_city##":"En avlägsen stad"
"##collapsed_building_text##":"En byggnad har rasat. Dåligt underhåll av stadens ingenjörer av orsakat detta."
"##day_longer_in_that_tent##":"En dag till i det tältet och jag hade exploderat"
"##nativeHut_info##":"En del lokalbefolkning bor här, de lever ett stillsamt enkelt liv. De vill bara bli lämnade ifred."
"##academy_info##":"En del ungdomar som går ut skolorna går vidare och studerar avancerad retorik och historia vid högskolan. Alla kulturella medborgare har en akademisk bakgrund."
"##wn_eygptian_soldier##":"En egyptisk soldat"
"##line_formation_text##":"En enkel formation, som ger fördelar åt försvarstrupper."
"##wn_etruscan_soldier##":"En etruskisk soldat"
"##pestilent_event_text##":"En farsot har drabbat staden. Bristen på sjukhus fordrar att dina prefekter desinfekterar de drabbade stadsdelarna."
"##enemy_army_threating_a_city##":"En fiendearmé som hotar en av rikets städer"
"##enemy_army_attack_city##":"En fiendes armé marserar i detta nu direkt mot dig stad. De har plundrat några städer i närheten, och de är beräknade att nå din stad detta år."
"##wn_gaul_soldier##":"En gallisk soldat"
"##blessing_of_mercury_title##":"En gåva från Merkurius"
"##blessing_of_neptune_title##":"En gåva från Neptunus"
"##goth_warrior##":"En gotisk soldat"
"##greek_soldier##":"En grekisk soldat"
"##egift_troupe_preforming_slaves##":"En grupp uppträdande slavar"
"##blessing_of_ceres_title##":"En gudagåva från Ceres"
"##spirit_of_mars_title##":"En gudagåva från Mars"
"##blessing_of_venus_title##":"En gudagåva från Venus"
"##egift_golden_chariot##":"En gyllene vagn"
"##wn_helveti_soldier##":"En helvetisk soldat"
"##hun_warrior##":"En hunnersoldat"
"##wn_iberian_soldier##":"En iberisk soldat"
"##judaean_warrior##":"En judéisk soldat"
"##wn_celt_soldier##":"En keltisk soldat"
"##emperror_legion_at_out_gates##":"En legion av kejsarens trupper står vid portarna"
"##small_fest_description##":"En liten festival hölls denna kväll. Alla är tacksamma över detta avbrott i vardagen."
"##macedonian_soldier##":"En makedonisk soldat"
"##defensive_formation_text##":"En mycket defensiv formation. Nästan omöjlig att penetreras av missiler."
"##nearby_building_negative_effect##":"En närliggande {0} har en försämrande effekt på efterfrågan till området. Försök att anlägga t ex trädgårdar, torg och statyer."
"##numidian_warrior##":"En numidisk soldat"
"##wt_pict_soldier##":"En piktisk soldat"
"##forum_information##":"En populär samlingsplats och eftertraktat samhällselement. Forum anställer även skatteindrivare och är livsviktiga för stadens skattkammare."
"##romechastener_attack_text##":"En romersk legion är inom sikte av staden. Detta är ett verkligen ett hot."
"##roman_city##":"En romersk stad"
"##samnite_soldier##":"En samnitisk soldat"
"##seleucid_soldier##":"En selucidisk soldat"
"##egift_soldier_from_pergamaum##":"En soldat från Pergamon"
"##egift_educated_slave##":"En utbildad slav"
"##wn_visigoth_soldier##":"En visigotisk soldat"
"##warehouse_no_workers##":"Endast minimibemanning. Kommer ej att sända eller ta emot varor"
"##formation_available_for_trained_troops##":"Endast tillgänglig för trupper som utbildats på militärhögskola."
"##wt_endeavor##":"Endeavor"
"##unit##":"Enhet"
"##employee##":"Enhet"
"##units##":"Enheter"
"##employees##":"Enheter"
"##tarentum_win_text##":"Etruskerna kommer inte att hota Tarentum igen. Bra gjort! Det är sällsynt med en ståthållare som finner rätt balans mellan stadsbyggnation och strid. Låt se om du kan göra om din bravad eller om det bara handlade om tur."
"##egift_gree_manuscript##":"Ett grekiskt manuskript"
"##lawless_area##":"Ett laglöst område. Människorna är vettskrämda."
"##fort_info##":"Ett romerskt fort rekryterar soldater från förläggningar. Lägga till en militärhögskola skulle ge trupper med bättre utbildning."
"##show##":"Evenemang"
"##god_exalted##":"Exalterad"
"##explosion##":"Explosion"
"##export##":"Export"
"##exports_over##":"Exportera vara över"
"##trade_btn_export_text##":"Exportera vara över"
"##extreme_fire_risk##":"Extrem brandrisk"
"##sldr_extremely_scared##":"Extremt rädd"
"##sldh_health_strongest##":"Extremt stark"
"##wn_eygptians##":"Eygptier"
"##wt_sheep##":"Får"
"##pestilence_event_text##":"Farsot"
"##high_bridge##":"Fartygsbro"
"##shipyard##":"Fartygsvarv"
"##export_btn_tooltip##":"Fastställ den kvantitet av dessa varor som du önskar behålla innan de exporteras"
"##setup_traderoute_to_import##":"Fastställ en handelsväg för att importera det"
"##wage_level_tip##":"Fastställ en lönenivå (ditt folk kommer att jämföra denna med lönerna i Rom)"
"##set_amount_to_donate##":"Fastställ summa att donera"
"##month_2_short##":"Feb"
"##festivals##":"Festivaler"
"##enemies_attack_title##":"Fiender attackerar staden"
"##barbarian_are_closing_city##":"Fiender närmar sig staden"
"##enemies_at_the_door##":"Fiender vid dina portar"
"##city_under_barbarian_attack##":"Fiendesoldaterna i stadens omgivning förbättrar inte din fredsställning!"
"##advchief_finance##":"Finanser"
"##finance_advisor##":"Stadens kapital"
"##finances##":"Finanser"
"##fish##":"Fisk"
"##fishing_boat##":"Fiskebåt"
"##fishing_wharf##":"Fiskehamn"
"##wharf##":"Fiskehamn"
"##fishing_waters##":"Fiskevatten"
"##healthadv_some_regions_need_doctors_2##":"Fler och fler människor vill ha bekväm tillgång till hälsovård. Anordna lokal tillgång till kliniker så att staden kan växa."
"##religionadv_need_basic_religion##":"Fler och fler medborgare kräver minst en gudstjänstplats i sitt bostadsområde, för att förbättra gudarnas uppfattning om dem."
"##healthadv_some_regions_need_barbers##":"Fler områden i staden kräver nu barberare. I takt med att din stad blir allt mer välbeställd kommer fler att ha tid till rakning och klippning!"
"##several_crimes_but_area_secure##":"Flera brott har rapporterats här nyligen, men på det hela taget har prefekterna situationen under kontroll"
"##cartPusher_average_life##":"Flytta kärror hela dagarna är knappast kul, men att leva här gör det möjligt."
"##bathlady_so_hungry##":"Folk har inte ätit på så länge att deras revben börjar sticka ut, vilket syns på badhuset."
"##money_stolen_title##":"Folket är arga"
"##citychart_census##":"Folkräkning"
"##fountain##":"Fontän"
"##for_second_year_broke_tribute##":"För andra året i rad har du inte betalat tribut till Rom. Detta håller på att bli ett stort problem för din framtida karriär."
"##no_room_for_citizens##":"för många"
"##too_close_to_enemy_troops##":"För nära fiendestyrkorna!"
"##prefecture_full_work##":"För närvarande är vår tjänstgöringslista full. Våra prefekter är alltid ute och patrullerar gatorna."
"##forum_full_work##":"För närvarande arbetar våra indrivare med maximal effektivitet, och de är alltid ute och kontrollerar att alla förfallna skatter betalas in till staden."
"##healthadv_not_need_health_service_now##":"För närvarande finns ingen efterfrågan på hälsovård eller sanitära inrättningar. I takt med att staden utvecklas, kommer dock befolkningen att kräva badhus och sjukhus, och senare även barberare!"
"##have_no_requests##":"För närvarande har du inga meddelanden att läsa. I takt med att din stad växer, eller om kejsaren begär varor av dig, kommer meddelanden att visas här"
"##engineering_post_full_work##":"För närvarande har vi inga driftavbrott Våra ingenjörer är alltid ute och inspekterar och reparerar skador på stadens byggnader."
"##entadv_small_city_not_need_entert##":"För tillfället har dina medborgare andra enklare behov, än underhållning att tänka på. Men i takt med att staden växer kommer de ha begär för något som minskar enformigheten i deras vardagsliv."
"##cursed_by_mars##":"Förbannad av Mars!"
"##prepare_to_festival##":"Förbereder den kommande festivalen"
"##smcurse_of_mercury_description##":"Förfärad över ditt bristande intresse för honom har Merkurius med andlig kraft avlägsnat en del varor från dina sädes- eller handelsmagasin."
"##wrath_of_ceres_description##":"Förgrummad över din brist av respekt mot Ceres, hon ger ditt folk en gräshopsplåga. Det kommer dröja innan dina grödor kan växa igen."
"##contaminted_water##":"Förorenat vatten"
"##last_year##":"Förra året"
"##lost_money_last_year##":"Förra året förlorade din stad pengar - detta minskade stadens välstånd."
"##emw_sell##":"Försäljningar"
"##landmerchant_say_about_store_goods##":"Försiktigt! Jag önskar att arbetarna skulle ta det lugnt när de lastar mina djur med de varor jag nyss har köpt."
"##granary_devastation_mode_text##":"Försöker att sända mat till annan plats"
"##warehouse_devastation_mode_text##":"Försöker sända gods till annan plats"
"##destroy_bridge##":"Förstör en bro"
"##destroy_fort##":"Förstör ett fort"
"##destroyed_building_title##":"Förstörd byggnad"
"##fort##":"Fort"
"##money_stolen_text##":"Fortfarande frustrerad, några invånare har börjat stjäla. De mer laglydiga invånarena har börjat prata om att flytta. Handla nu för att förbättra humöret på dem."
"##blessing_of_ceres_description##":"Förtjust över den uppmärksamhet som din stad visar henne förbättrar Ceres fruktbarheten hos din växande gröda."
"##blessing_of_mercury_description##":"Förtjust över din hängivenhet har Merkurius upptäckt bortglömda produkter i ett av stadens sädesmagasin."
"##delighted##":"Förtjusta"
"##continue##":"Fortsätt"
"##mainmenu_continueplay##":"Fortsätt"
"##plname_continue##":"Fortsätt"
"##continue_2_years##":"Fortsätt att styra i 2 år till."
"##continue_5_years##":"Fortsätt i 5 år till."
"##forum##":"Forum"
"##qty_stacked_in_city_warehouse##":"förvaras i stadens handelsmagasin"
"##message_from_centurion##":"Från legion's centurion..."
"##senatepp_peace_rating##":"Fred"
"##wndrt_peace##":"Fredsställning"
"##peace_rating_text##":"Fredsställningen blir bättre för varje år utan upplopp eller invasioner som skadar egendom i städerna."
"##egift_lavish##":"Frikostig:"
"##fruit##":"Frukt"
"##fig_farm_info##":"Frukt är en viktig del av den balanserad diet som ditt folk behöver för hälsa och glädje. I sädesmagasinen lagras frukt för lokal konsumtion, och i handelsmagasinen förvaras överskottet för export."
"##fig_farm##":"Fruktodling"
"##granary_info##":"Fulla sädesmagasin är livsviktiga för att hålla folkets magar fyllda och för att attrahera nya medborgare. Ett sädesmagasin kan lagra säd, kött, grönsaker och frukt."
"##fullscreen_on##":"Fullskärm"
"##need_barracks_for_work##":"Fungerande förläggning krävs för att ta emot soldater"
"##working_industry##":"fungerande industri i staden"
"##working_industries##":"fungerande industrier i staden"
"##empbutton_low_work##":"Fungerar dåligt. Tilldela fler människor till vår sektor"
"##factory_need_more_workers##":"Fungerar knappt. Tilldela fler människor till vår sektor"
"##empbutton_simple_work##":"Fungerar, men fler arbetare skulle kunna tilldelas oss"
"##goto##":"Gå till"
"##empire_map##":"Gå till imperiet"
"##goto_empire_map##":"Gå till kartan över imperiet"
"##disasterBtnTooltip##":"Gå till problemområde."
"##wn_gaul##":"Galler"
"##egift_gaulish_bodyguards##":"Galliska livvakter"
"##give_money##":"Ge pengar"
"##send_money_to_city##":"Ge pengar till staden"
"##send_to_city##":"Ge till staden"
"##overall_people_are_coming_city##":"Generellt sett, kommer folket till din stad, eller vill de komma."
"##overall_people_are_leaving_city##":"Generellt sett, lämnar folket din stad."
"##egift_generous##":"Generös:"
"##egift_gepards_and_giraffes##":"Geparder och giraffer"
"##may_collect_about##":"ger en avkastning på"
"##blessing_of_neptune_description##":"Glad över ditt växande intresse för honom garanterar Neptunus alla dina sjöfarande handelsmän lugna seglatser under resten av året. De kommer att betala dig dubbelt under den tiden."
"##god_happy##":"Glada"
"##wt_gladiator##":"Gladiator"
"##gladiator_bouts_runs_for_another##":"Gladiatorkampen pågår ytterligare"
"##gladiator_pit##":"Gladiatorskola"
"##gladiatorSchool##":"Gladiatorskola"
"##sldh_health_sparse##":"Gles"
"##empireBtnTooltip##":"Global karta"
"##gmenu_shortkeys##":"Globala kortkommandon"
"##no_dock_for_sea_trade_routes##":"GLÖM INTE! Denna nya handelsrutt över havet kräver byggnation av en handelshamn innan några fartyg kan anlända."
"##marketBuyer_good_life##":"God dag, medborgare. Är det inte en härlig stad?"
"##minimizeBtnTooltip##":"Göm panel"
"##hide_bigpanel##":"Göm sidopanelen, och utöka spelvyn"
"##trade_btn_notrade_text##":"Gör ej affärer"
"##wn_goth##":"Gother"
"##graphics##":"GRAFIK:"
"##grass##":"Gräs"
"##congratulations##":"Gratulerar"
"##tutorial_win_text##":"Gratulerar! Du har förstått grunderna på ett nöjsamt sätt. För att på bästa sätt fortsätta din utbildning, har jag ännu ett lindrigt uppdrag åt dig. Mot Brundisium!"
"##ive_asked_senate_proclaim_you_a_god##":"Gratulerar! Du har uppnått de högsta poängställningar som någonsin åstadkommits av Roms ståthållare. Jag är stolt över att få lämna över till dig. Jag kungör att du må krönas till kejsare och härskare över hela imperiet. Äntligen kan jag dra mig tillbaka till min villa på ön, som en vanlig medborgare igen. Må ditt namn..."
"##wn_graeci##":"Greker"
"##gatehouse##":"Grindstuga"
"##vegetable##":"Grönsaker"
"##vegetable_farm_info##":"Grönsaker är en viktig del av den balanserad diet som ditt folk behöver för hälsa och glädje. I sädesmagasinen lagras grönsaker för lokal konsumtion, och i handelsmagasinen förvaras överskottet för export."
"##vegetable_farm##":"Grönsaksodling"
"##gods_unhappy_title##":"Gudar är missnöjda"
"##city_opts_god_off##":"Gudar: Av"
"##city_opts_god_on##":"Gudar: På"
"##rladv_mood##":"Gudarna är"
"##lionTamer_gods_angry##":"Gudarna är så rasande att det påverkar mitt Lejon! Han är rytande arg!"
"##gods_wrathful_title##":"Gudarna är vreda"
"##god_neptune_short##":"Guden Neptune..."
"##favor##":"Gynna"
"##senatepp_favour_rating##":"Gynna"
"##wndrt_favour##":"Gynna"
"##advchief_health##":"Hälsa"
"##health##":"Hälsa"
"##healthAll##":"Hälsa"
"##ovrm_health##":"Hälsa"
"##healthBtnTooltip##":"Hälsa"
"##wt_docker##":"Hamnarbetare"
"##dockers_taking_our_goods##":"Hamnarbetarna för våra varor till lagerlokalen nu."
"##dock_info##":"Handelsskepp från hela riket lägger till här för att leverera importvaror och hämta exportvaror. Du kan inte bedriva sjöhandel utan en handelshamn."
"##stacking##":"Hamstrar"
"##stacking_resource##":"Hamstrar vara"
"##deliver##":"Hämta varor"
"##ovrm_commerce##":"Handel"
"##mercury_desc##":"Handel"
"##trade##":"Handel"
"##comerceBtnTooltip##":"Handel"
"##commerce##":"Handel"
"##dock##":"Handelshamn"
"##warehouse##":"Handelsmagasin"
"##warehouses##":"Handelsmagasin"
"##small_mercury_temple_info##":"Handelsmännen dyrkar Merkurius för att skydda sina varor. Om Merkurius vrede väcks sätts allas vinst på spel."
"##trade_advisor##":"Handelsrådgivare"
"##trade_ship_from##":"Handelsskepp från"
"##no_working_dock##":"Handelsskepp från hela riket lägger till här för att leverera importvaror och hämta exportvaror. Du kan inte bedriva sjöhandel utan en handelshamn."
"##lionTamer_average_life##":"Här är lite utländskt kött åt dig, Leo."
"##imperial_reminder_text##":"Har du glömt bort min senaste förfrågan? Jag börjar tappa tålamodet."
"##taxCollector_high_tax##":"Har du sett skatterna här? Medborgare, det är inte rätt."
"##pottery_workshop_info##":"Här formar krukmakare lera till kärl som medborgarna använder till förvaring. Handla med krukor, eller låt dina marknader distribuera dem så att människorna kan bygga bättre hus."
"##patrician_average_life##":"Här i min bekväma villa anser jag livet i staden vara mycket bra."
"##waiting_for_free_dock##":"Har kastat ankar, i väntan på ledig kajplats"
"##oil_workshop_info##":"Här pressas olja från oliver, som plebejerna behöver för matlagning och för belysningen i sin Insulae. Överskottsoljan kan bli lönsam handel."
"##game_speed_options##":"Hastighetsinställningar"
"##speed_settings##":"Hastighetsinställningar"
"##neptune_desc##":"Havet"
"##patrician_so_hungry##":"Hell! Vad tjänar rikedom till om det inte finns mat att köpa?"
"##wt_homeless##":"Hemlös"
"##prefect_fight_fire##":"Hettan från elden är otroligt stark."
"##lgn_stallion##":"Hingstarna"
"##hippodrome##":"Hippodrom"
"##ovrm_hippodrome##":"Hippodrom"
"##hippodromes##":"Hippodromer"
"##valencia_win_text##":"Hispaniens nya huvudstad är precis vad vi behöver för att knyta den avlägsna provinsen tätare till Rom. Genom att krossa etruskerna så totalt försvinner det sista hotet i väst."
"##citychart_population##":"Historia"
"##no_tax_in_this_year##":"Hittills i år har ingen skatt betalats från detta hus"
"##gmenu_help##":"Hjälp"
"##help##":"Hjälp"
"##scholar_gods_angry##":"Hjälp! Gudarna är vreda. De kommer att straffa oss."
"##lgn_heroes##":"Hjältarna"
"##migration_broke_workless##":"Hög arbetslöshet i din stad bromsar din välståndsställning."
"##migration_lack_crime##":"Hög brottslighet skrämmer lokalbefolkningen."
"##migration_lack_tax##":"Höga skatter är ett problem"
"##migration_middle_lack_tax##":"Höga skatter förhindrar immigration"
"##migration_broke_tax##":"Höga skatter gör att vissa människor undviker din stad"
"##press_escape_to_exit##":"Högerklicka för att avsluta"
"##right_click_to_exit##":"Högerklicka för att avsluta"
"##colleges##":"Högskolor"
"##mainmenu_dlc_main##":"Hur man bygger Rom"
"##romeGuard_so_hungry##":"Hur ska en soldat kunna slåss utan mat?"
"##houseBtnTooltip##":"Hus"
"##lgn_hydras##":"Hydrorna"
"##library_no_workers##":"Hyllorna i detta bibliotek är tomma, och värdelösa för lokalsamhället."
"##work##":"I bruk"
"##entertainment_need_for_upgrade##":"I delar av staden klagar man över frånvaron av fritidsanläggningar. Byggnation av fler platser för underhållning skulle hjälpa utvecklingen i de fattigare områdena."
"##romeGuard_high_workless##":"I dessa tider av arbetslöshet tackar jag gudarna att jag har jobb."
"##students##":"i högskoleålder."
"##your_salary_frowned_senate##":"I Rom ser man ner på din fräckhet att betala dig själv en lön som är högre än din rang."
"##scholars##":"i skolålder"
"##senate_save##":"i stadskassan"
"##wt_immigrant##":"Immigrant"
"##emperor##":"Imperiet"
"##RomeChastenerArmy_troops_at_our_gates##":"Imperiets trupper står vid stadsportarna"
"##import_fn##":"Importer"
"##import##":"Importerar"
"##trade_btn_import_text##":"Importerar"
"##industry_disabled##":"Industri är AV"
"##industry_enabled##":"Industri är PÅ"
"##wt_indigene##":"Inföding"
"##wn_indigene##":"Infödingar"
"##native_hut##":"Infödingshydda"
"##colloseum_haveno_animal_bouts##":"Inga djurkamper för närvarande"
"##no_industries_in_city##":"Inga industrier i staden"
"##hippodrome_haveno_races##":"Inga kapplöpningar för närvarande"
"##no_people_in_city##":"Inga människor i staden!"
"##no_people_in_this_locality##":"Inga människor på denna plats."
"##not_need_education##":"Inga medborgare kräver ännu utbildningsmöjligheter. Men när staden börjar växa kommer människor att förvänta sig skolor och högskolor, och senare även bibliotek."
"##no_citizens_desire_live_here##":"Inga medborgare vill bo här"
"##srcw_no_messages##":"Inga nya meddelanden"
"##colloseum_haveno_gladiator_bouts##":"Ingen aktuell gladiatorkamp"
"##no_fire_risk##":"Ingen brandrisk"
"##none_crime_risk##":"Ingen brottslighet i sikte här."
"##freehouse_text##":"Ingen har så mycket som satt upp ett tält här ännu, fast immigranter kommer säkert att anlända inom kort om staden har tillgång till livsmedel och arbeten."
"##freehouse_text_noroad##":"Ingen kommer att skapa sig ett hem här eftersom det ligger för långt från närmaste väg. Om ingen väg byggs snart kommer detta område att återgå till öppet landskap."
"##no_food_stored_last_month##":"INGEN MAT lagrad förra månaden!"
"##no_priority##":"Ingen prioritet"
"##none_damage_risk##":"Ingen risk för kollaps"
"##engineer##":"Ingenjör"
"##wt_engineer##":"Ingenjör"
"##engineering_post_info##":"Ingenjörer är mycket respekterade yrkesmän, och det är alltid stor efterfrågan på deras tjänster. Konstant underhåll förhindrar att byggnaderna faller samman."
"##engineering_structures##":"Ingenjörsbyggnader"
"##engineer_salary##":"Ingenjörslön på"
"##engineering_post##":"Ingenjörspostering"
"##ovrm_simple##":"Ingenting"
"##landmerchart_noany_trade2##":"Inget att byteshandla med här, passerar bara"
"##hippodrome_no_workers##":"Inget rör sig i hippodromen. Utan arbetare ger den ingen underhållning åt lokalsamhället."
"##missionaryPost##":"Inhemsk mission"
"##native_center##":"Inhemskt centrum"
"##taxes##":"Inkasserade skatter"
"##debet##":"Inkomst"
"##emw_buy##":"Inköp"
"##options##":"Inställning"
"##warehouse_orders##":"Instruktioner handelsmagasin"
"##granary_orders##":"Instruktioner sädesmagasin"
"##pop##":"Inv"
"##overall_city_population_static##":"Invånarantalet i din stad är i stort sett statiskt."
"##occupants##":"invånare"
"##lowgrade_housing_want_better_conditions##":"Invånarna i dåliga bostäder vill ha bättre villkor"
"##city_zoominv_off##":"Inverterad zoom: Av"
"##city_zoominv_on##":"Inverterad zoom: På"
"##yes##":"Ja"
"##taxСollector_much_tax##":"Jag älskar att driva in skatt från rika hus som dessa."
"##landmerchant_good_deals##":"Jag älskar att komma hit. Affärerna går mycket bra."
"##merchant_little_busy_now##":"Jag är lite upptagen just nu."
"##emperor_wrath_by_debt_text##":"Jag är mycket missnöjd. Trots alla pengar jag har investerat i din stad och senatens generösa krediter, har du svikit mig. Din stad har inte betalat tillbaka sina lån. Mitt förtroende för dig var missriktat och jag tvingas nu finna en annan ståthållare i ditt ställe. Du kanske passar bättre i den nya position jag har i åtanke för dig..."
"##immigrant_where_my_home##":"Jag är ny i staden. Vet du var man kan få tag i en bostad?"
"##prefect_gods_angry##":"Jag är rädd för att gudarna kommer att förbanna staden."
"##wt_missioner_normal_life##":"Jag är så glad att vara romare. Du skulle se vad dessa barbarer håller på med i sina hyddor!"
"##gladiator_so_hungry##":"Jag är så hungrig att jag kan äta ett lejon!"
"##recruter_low_entertainment##":"Jag arbetar hårt och jag vill roa mig ofta. Men det går inte här. Det finns inget att göra!"
"##engineer_building_allok##":"Jag behövs knappast. Dessa byggnader är i utmärkt skick."
"##legionary_low_salary##":"Jag får inte tillräckligt bra betalt för att slåss!"
"##rome_need_some_money##":"Jag ger dig härmed förmånen att tillhandahålla ytterligare medel för det goda i Rom. Skicka dem snart, och jag kommer att överväga att konstruera en staty i din ära."
"##marketBuyer_need_workers##":"Jag har aldrig sett så många byggnader som behöver fler arbetare."
"##emigrant_thrown_from_house##":"Jag har blivit utkastad från mitt hem!"
"##emigrant_no_work_for_me##":"Jag har fått nog av detta ställe. Det finns inget arbete här."
"##lion_pit_bad_work##":"Jag har ingen personal utöver mig själv. Jag kan inte arbeta under dessa förhållanden! Som bäst kan jag leverera ett lejon på tre månader."
"##gladiator_pit_bad_work##":"Jag har ingen personal utöver mig själv. Jag kan inte arbeta under dessa förhållanden! Som bäst kan jag utbilda en gladiator var tredje månad."
"##emigrant_no_home##":"Jag har ingenstans att bo."
"##merchant_notbad_city##":"Jag har kappkört i många värre städer än den här."
"##romeGuard_good_live##":"Jag må vara en simpel soldat, men även jag kan se vilken storslagen stad detta är."
"##taxCollector_high_workless##":"Jag ogillar det här stället. Arbetslösheten är för hög."
"##marketBuyer_find_goods##":"Jag ska hämta nya varor."
"##taxCollector_low_entertainment##":"Jag skulle inte ha nåt emot att pressa folk på denarer hela dagarna om det bara fanns mer att göra på kvällarna!"
"##legionary_average_life##":"Jag slåss intill döden! Staden är trygg så länge jag lever!"
"##landmerchant_noany_trade##":"Jag vet inte varför jag tar den här handelsvägen. De köper ingenting och de har inget de vill sälja till mig."
"##merchant_wait_for_deal##":"Jag vill gärna göra affärer här. Jag älskar att göra en bra affär."
"##month_1_short##":"Jan"
"##iron##":"Järn"
"##earthquake_title##":"Jordbävning"
"##ceres_desc##":"Jordbruk"
"##trouble_farm_was_blighted_by_locust##":"Jordbrukets marker har skadats av gräshoppssvärmarna, återhämtningen kommer att ta tid."
"##wn_judaean##":"Judeér"
"##month_7_short##":"Juli"
"##month_6_short##":"Juni"
"##recruter_so_hungry##":"Kan du avvara lite bröd? Jag har inte ätit på så länge."
"##water_info##":"Kan inte forceras, men broar kan byggas på vissa platser. Vatten är en vital handelslänk till resten av imperiet via handelshamnar. Lertag måste byggas nära vatten."
"##unable_fullfill_request##":"Kan inte fullgöra begäran"
"##lgn_rabbits##":"Kaninerna"
"##current_races_runs_for_another##":"Kapplöpningar pågår ytterligare"
"##venus_desc##":"Kärlek"
"##wn_carthaginians##":"Karthager"
"##funds_tooltip##":"Kassa"
"##fort_javelin##":"Kastspjut"
"##earthquake_text##":"Katastrof! Till och med gudarna är chockade. En jordbävning som sväljer allt i sin väg. Hoppas det går bra, reparera alla skador när det slutar."
"##lutetia_win_text##":"Kejsar Augustus måste ha anat ditt styre när han förutspådde vår seger över gallerna. Din framgång vid Lutetia räcker långt när det gäller att krossa deras upprorsanda."
"##emperor_favour_04##":"Kejsaren är arg på dig."
"##emperor_favour_16##":"Kejsaren är entusiastisk över vad du gjort."
"##emperor_favour_17##":"Kejsaren är extremt entusiastisk över vad du gjort."
"##emperor_favour_05##":"Kejsaren är extremt missnöjd med dig."
"##emperor_favour_10##":"Kejsaren är fundersam vad gäller dig."
"##emperor_favour_19##":"Kejsaren är mer än tillfreds med vad du gjort."
"##emperor_favour_07##":"Kejsaren är missnöjd med dig."
"##emperor_favour_03##":"Kejsaren är mycket arg på dig."
"##emperor_favour_14##":"Kejsaren är mycket entusiastisk över vad du gjort."
"##emperor_favour_06##":"Kejsaren är mycket missnöjd med dig."
"##emperor_favour_13##":"Kejsaren är mycket nöjd med vad du gjort."
"##emperor_favour_08##":"Kejsaren är något missnöjd med dig."
"##emperor_favour_15##":"Kejsaren är nöjd med vad du gjort."
"##emperor_favour_00##":"Kejsaren är rasande på dig."
"##emperor_favour_01##":"Kejsaren är så otroligt arg att han talar om att landsförvisa dig."
"##emperor_favour_20##":"Kejsaren är så otroligt nöjd att han talar om att utnämna dig till sin arvinge."
"##emperor_favour_12##":"Kejsaren är tillfreds med dig."
"##emperor_favour_09##":"Kejsaren är tveksam vad gäller dig."
"##emperor_favour_18##":"Kejsaren är utom sig av glädje över vad du gjort."
"##emperor_favour_02##":"Kejsaren är vansinnigt arg på dig."
"##emperor_limit_houseupgrade##":"Kejsaren har begränsat uppgraderingar av husen i denna stad"
"##emperor_favour_11##":"Kejsaren tror du kan bevisa dig värdefull ."
"##wn_celts##":"Kelter"
"##wt_surgeon##":"Kirurg"
"##emperor_request_money##":"Kjesare efterfrågar pengar"
"##emperor_request##":"Kjesare efterfrågar varor"
"##city_still_in_debt_text##":"Kjesaren är rasande på dig för att du fortfarande är skylldig Rom pengar. Han ger dig 12 månader till att betala skulden. Annars kommer du straffas ordentligt."
"##its_very_peacefull_province##":"Kjesaren har aldrig förut skådat en sådan fridfull stad förut!"
"##emperor_anger##":"Kjesarens ilska"
"##rome_gratitude_request_title##":"Kjesarens tacksamhet."
"##advemp_emperor_favour##":"Kjeserlig förmån"
"##imperial_reminder##":"Kjeserlig påminnelse"
"##legion_formation_tooltip##":"Klicka här för att ändra legionens formation"
"##restart_mission_tip##":"Klicka här för att återuppbygga denna provins"
"##give_money_tip##":"Klicka här för att donera pengar till staden"
"##set_mayor_salary##":"Klicka här för att fastställa din personliga lön"
"##empbutton_tooltip##":"Klicka här för att fastställa en prioritet för denna arbetskraftskategori"
"##go_to_problem##":"Klicka här för att gå till detta problemområde"
"##click_here_that_stacking##":"Klicka här för att hamstra"
"##request_btn_tooltip##":"Klicka här för att sända iväg begäran"
"##click_here_that_use_it##":"Klicka här för att stänga av hamstring"
"##click_here_to_talk_person##":"Klicka här för att tala med denna person"
"##wndrt_peace_tooltip##":"Klicka här för information om din fredsställning"
"##wndrt_favor_tooltip##":"Klicka här för information om din popularitetsställning"
"##wndrt_prosperity_tooltip##":"Klicka här för information om din välståndsställning"
"##minimap_tooltip##":"Klicka på denna översiktskarta för att flytta till avlägsna delar av din stad"
"##click_on_city_for_info##":"Tryck på stad för information"
"##click_item_for_start_trade##":"Klicka på en vara"
"##priority_button_tolltip##":"Klicka på ett nummer för att fastställa prioritetsnivå. Alla övriga uppgifter kommer att omjusteras"
"##clinic##":"Klinik"
"##ovrm_clinic##":"Kliniker"
"##clinics##":"Kliniker"
"##rock_caption##":"Klippor"
"##rock_text##":"Klipporna kan inte forceras eller röjas undan. Marmor- och malmbrott fungerar bara om de uppförs nära klippor."
"##collapsed_building_title##":"Kollapsad byggnad"
"##column_info##":"Kolonnformation"
"##consul##":"Konsul"
"##consul_salary##":"Konsulslön på"
"##buy_price##":"Köparna betalar"
"##trade_caravan_from##":"Köpmannakaravan från"
"##emw_bought##":"Köpt"
"##marketKid_say_2##":"Korgen tar kål på mig. Jag bryr mig inte om vem som behöver maten, det borde finnas en lag mot barnarbete."
"##cost##":"Kostnad"
"##cost_2_open##":"Kostnad att öppna"
"##costs##":"kostnader"
"##meat##":"Kött"
"##demand##":"Krav"
"##demands_3_religion##":"Krav på tillgång till en tredje religion"
"##rioter_rampaging_accross_city##":"Kravaller i staden. De förstör och tar allt de kommer över."
"##need_access_to_full_reservoir##":"Kräver tillgång till en full reservoar för att fungera"
"##need_population##":"krävs)"
"##out_of_credit##":"Kredit saknas!"
"##mars_desc##":"Krig"
"##migration_war_deterring##":"Krig avskräcker immigranter!!"
"##pottery_workshop##":"Krukmakeri"
"##pottery##":"Krukor"
"##senatepp_clt_rating##":"Kultur"
"##wndrt_culture##":"Kultur"
"##coast_caption##":"Kuster"
"##quaestor_salary##":"Kvestorslön på"
"##load_this_game##":"Ladda"
"##start_this_map##":"Starta denna karta"
"##mainmenu_loadcampaign##":"Ladda kampanj"
"##mainmenu_playmission##":"Ladda scenario"
"##mainmenu_load##":"Ladda spel"
"##mainmenu_loadgame##":"Ladda spel"
"##initialize_animations##":"Laddar animationer"
"##initialize_walkers##":"Laddar fotgängarinställningar"
"##initialize_house_specification##":"Laddar husdata"
"##initialize_constructions##":"Laddar konstruktionsinställningar"
"##initialize_names##":"Laddar medborgarnamnen"
"##initialize_religion##":"Laddar religioninställningar"
"##loading_offsets##":"Laddar texturer"
"##loading_resources##":"Laddar tillgångar"
"##low_bridge##":"Låg bro"
"##low_wage_lack_migration##":"Låga löner är ett problem"
"##low_wage_broke_migration##":"Låga löner minskar immigrationen till din stad"
"##merchant_just_unloading_my_goods##":"Lagerlokalen lastar just av varor från mina djur."
"##grape_factory_stock##":"Lagrade druvor,"
"##olive_factory_stock##":"Lagrade oliver,"
"##units_in_stock##":"Lagrar"
"##iron_factory_stock##":"Lagrat järn,"
"##timber_factory_stock##":"Lagrat virke,"
"##clinic_info##":"Läkares förbättrar medborgarnas hälsa genom sina hembesök i de stadsdelar som ingår i deras runda. Blomstrande områden vill ha en klinik."
"##leave_empire?##":"Lämna det Romerska Riket?"
"##donationwnd_exit_tip##":"Lämna donationsskärmen"
"##exit_salary_window##":"Lämna löneskärmen"
"##land_route##":"Landväg"
"##farm##":"Lantbruk"
"##wt_teacher##":"Lärare"
"##free##":"ledig"
"##freehouse_caption##":"Ledig tomt"
"##wt_legioanry##":"Legionär"
"##fort_legionaries##":"Legionärfort"
"##legion_morale_is_too_low##":"Legionens stridsmoral är för dålig för att kunna svara!"
"##legions##":"Legioner"
"##romechastener_attack_title##":"Legioner anfaller"
"##lgn_lions##":"Lejonen."
"##lion_pit##":"Lejonhus"
"##lionsNusery##":"Lejonhus"
"##wt_lion_tamer##":"Lejontämjare"
"##lionTamer_low_entertainment##":"Leo och jag slåss dygnet runt och ändå har folk tråkigt. Det finns helt enkelt inte tillräckligt med artister här."
"##docked_buying_selling_goods##":"Ligger vid kaj, köper och säljer varor"
"##god_indifferent##":"Likgiltiga"
"##lindum_title##":"Lindum: en extremt farlig provins"
"##line_formation_title##":"Linjeformation"
"##low_fire_risk##":"Liten brandrisk"
"##small_festival##":"Liten festival"
"##small_domus##":"Liten Insulae"
"##small_shack##":"Liten koja"
"##low_damage_risk##":"Liten risk att kollapsa"
"##status_small##":"Liten staty"
"##small_villa##":"Liten villa"
"##small##":"Litet"
"##small_hut##":"Litet hus"
"##small_palace##":"Litet palats"
"##small_hovel##":"Litet skjul"
"##small_tent##":"Litet tält"
"##library_info##":"Litterära arbeten från hela riket förvaras här på grekiska och latin. Lärda män insisterar att biblioteken är avgörande för en viktig stad."
"##sldr_terrified##":"Livrädd"
"##have_food_for##":"Livsmedelsförråd för"
"##game_sound_options##":"Ljudalternativ"
"##gmsndwnd_ambient_sound##":"Ljudeffekter"
"##mainmenu_sound##":"Ljudinställningar"
"##sound_settings##":"Ljudinställningar"
"##localization##":"LOKALISERING:"
"##londinium_title##":"Londinium: une province pacifique"
"##advemployer_panel_salary##":"Löner"
"##wages##":"Löner"
"##lugdunum_title##":"Lugdunum: une province pacifique"
"##lutetia_title##":"Lutetia: une province dangereuse"
"##luxury_palace##":"Lyxpalats"
"##warehouseman##":"Magasinsman"
"##month_5_short##":"Maj"
"##mission_wnd_targets_title##":"Mål"
"##iron_mine##":"Malmbrott"
"##iron_mine_collapse##":"Malmbrott kollapsar"
"##months_until_defeat##":"Månader till nederlag"
"##months_until_victory##":"Månader till seger"
"##months##":"Människor"
"##months_to_comply##":"Människor"
"##people_leave_city_low_wage##":"Människor beger sig av på jakt efter högre löner"
"##road_paved_text##":"Människor föredrar torg!"
"##migration_peoples_arrived_in_city##":"Människor immigrerar till staden"
"##people_leave_city_some##":"Människor lämnar staden"
"##people_leave_city_insane_tax##":"Människor lämnar staden på grund av dina höga skatter"
"##more_4_month_from_festival##":"Människor talar fortfarande varmt om din senaste festival."
"##sentiment_people_love_you##":"Människorna älskar dig"
"##sentiment_people_angry_you##":"Människorna är arga på dig"
"##sentiment_people_extr_pleased_you##":"Människorna är extremt nöjda med dig"
"##sentiment_people_annoyed_you##":"Människorna är irriterade på dig"
"##sentiment_people_indiffirent_you##":"Människorna är likgiltiga inför dig"
"##sentiment_people_veryangry_you##":"Människorna är mycket arga på dig"
"##sentiment_people_verypleased_you##":"Människorna är mycket nöjda med dig"
"##sentiment_people_veryupset_you##":"Människorna är mycket upprörda över dig"
"##sentiment_people_pleased_you##":"Människorna är nöjda med dig"
"##sentiment_people_upset_you##":"Människorna är upprörda över dig"
"##sentiment_people_idolize_you##":"Människorna avgudar dig, som en gud"
"##fountain_info##":"Människorna hämtar allt vatten som de behöver från fontäner, som måste förses med vatten via ledningar från en reservoar. Fontäner är den källa till vatten som folket föredrar."
"##more_16_month_from_festival##":"Människorna kommer inte längre ihåg den sista festivalen som hölls i staden."
"##month_3_short##":"Mar"
"##market##":"Marknad"
"##marketLady_no_food_on_market##":"Marknaden har slut på livsmedel, så jag är på väg hem."
"##wt_marketBuyer##":"Marknadsbesökare"
"##wt_marketLady##":"Marknadshandlare"
"##ovrm_market##":"Marknadstillgång"
"##marble##":"Marmor"
"##quarry##":"Marmorbrott"
"##god_mars_short##":"Mars"
"##smallcurse_of_mars_title##":"Mars är upprörd"
"##wrath_of_mars_text##":"Mars börjar bli arg på dig. Le om du vågar. Fastän du inte har några millitärastyrkor idag. Mars blir inte så lätt förolämpad. Va vaksam!"
"##smallcurse_of_mars_description##":"Mars ogillar din brist på vördnad och sporrar ett antal missnöjda invånare att revoltera."
"##smallcurse_of_mars_text##":"Mars, soldaternas beskyddare och segerförlänare, är missnöjd. Dina soldater fruktar att de kommer att förlora ett stort slag om han inte blidkas."
"##wrath_of_mars_title##":"Mars vrede"
"##smallcurse_of_mars_failed_title##":"Mars vrede"
"##small_mars_temple##":"Marstempel"
"##massilia_title##":"Massilia: une province pacifique"
"##tower_need_wall_for_patrol##":"Måste finnas intill en mur för att sända ut en patrull"
"##ovrm_food##":"Mat"
"##advchief_food_consumption##":"Matförbrukning"
"##wharf_full_work##":"Med fullt antal anställda lassar och lossar vi med maximal hastighet."
"##barracks_have_weapons_bad_workers##":"Med minimipersonal utbildar vi nya soldater mycket långsamt trots att vi har de vapen som krävs för att utbilda alla typer av soldater."
"##shipyard_info##":"Med några vagnslaster timmer och tillräckligt med arbetare bygger fartygsvarvet fiskebåtar till stadens fiskehamnar."
"##olive_farm_bad_work##":"Med nästan inga anställda här, de flesta olivträd saknar oliver."
"##oil_workshop_bad_work##":"Med nästan inga anställda i olivodlingen, har produktionen avtagit. Det kommer produceras mycket lite olivolja det kommande året."
"##fruit_farm_slow_work##":"Med nästan inga anställda vid dem här fruktodlingen, kommer det ta evigheter att få någon frukt här."
"##quarry_bad_work##":"Med nästan inga anställda vid det här stenbrottet. Det kommer inte att produceras mycket marmor det kommande året."
"##iron_mine_bad_work##":"Med nästan inga gruvarbetare här, står nästan produktionen helt still. Det kommer inte produceras mycket järn det kommande året."
"##furniture_workshop_bad_work##":"Med nästan inga snickare i verkstan, står produktionen nästan stilla. Det kommer inte att produceras mycket möbler under det kommande året."
"##wine_workshop_bad_work##":"Med så få anställda står produktionen nästan still. Det kommer att produceras mycket lite vin under det kommande året."
"##weapons_workshop_bad_work##":"Med så få anställda står produktionen nästan still. Det kommer inte att produceras många vapen under det kommande året."
"##pottery_workshop_bad_work##":"Med så få anställda vid krukmakeriet står produktionen nästan stilla. Det kommer inte att produceras mycket krukor under det kommande året."
"##citizen##":"Medborgare"
"##etertadv_as_city_grow_you_need_more_entert##":"Medborgare som söker tidsfördriv har allt vad de behöver. Men i takt med att staden växer måste du förse dem med mer storslagen form av underhållning."
"##well_info##":"Medborgare utan tillgång till fontän kan ta vatten från brunnar, men stadsdelar med brunnsvatten är inga trevliga platser att bo på."
"##recruter_need_workers##":"Medborgare! Denna stad behöver fler arbetare."
"##gladiator_perfect_life##":"Medborgare! Jag har kämpat i många städer och den här är en av de bästa."
"##patrician_gods_angry##":"Medborgare! Situationen är hotfull. Gudarna är vreda."
"##citizens_here_are_bored_for_chariot_races##":"Medborgarna är uttråkade. Trots hästkapplöpningarna finns det inte tillräckligt med underhållning här."
"##gods_wrathful_text##":"Medborgarna fruktar att minst en av gudarna hyser vrede mot staden. De bönfaller dig att bygga fler tempel för att blidka dem."
"##religionadv_need_second_religion##":"Medborgarna i vissa områden vill ha tillgång till en annan religion nära hemmet. Bristen på religioner hindrar stadens utveckling i vissa områden."
"##citizens_grumble_lack_festivals_held##":"Medborgarna klagar över bristen på festivaler i din stad."
"##advchief_some_need_education##":"Medborgarna kräver mer utbildning"
"##citizens_enjoy_drama_and_comedy##":"Medborgarna njuter av drama och komedi enligt den grekiska traditionen."
"##citizens_like_chariot_races##":"Medborgarna vet inget bättre än vagnkapplöpningar."
"##message##":"Meddelande"
"##messages##":"Meddelanden"
"##messageBtnTooltip##":"Meddelanden från dina skrivare"
"##scribe_messages_title##":"Meddelanden från dina skrivare"
"##middle_insula##":"Medelstor Insulae"
"##statue_middle##":"Medelstor staty"
"##middle_villa##":"Medelstor villa"
"##middle_palace##":"Medelstort palats"
"##mediolanum_title##":"Mediolanum: province très dangereux"
"##mercury##":"Mercury"
"##smallcurse_of_mercury_failed_title##":"Mercury is upprörd"
"##smallcurse_of_mercury_title##":"Mercury is upprörd"
"##wrath_of_mercury_description##":"Mercury kokar av ilska. Brinnande stenar faller från himlen, som förstör byggnader och dess innehåll!"
"##wrath_of_mercury_title##":"Mercury vrede"
"##smcurse_of_mercury_title##":"Merkurius är upprörd"
"##smallcurse_of_mercury_description##":"Merkurius, gudarnas budbärare och handelsmännens beskyddare, är missnöjd. Dina handelsmän fruktar att hans beskydd viker."
"##small_mercury_temple##":"Merkuriustempel"
"##month##":"Mes"
"##month_to_comply##":"Mes"
"##miletus_title##":"Milet: province largement pacifique"
"##legion##":"Militär"
"##militaryAcademy##":"Militärhögskola"
"##more_8_month_from_festival##":"Minnet av den tidigare festivalen håller på att blekna."
"##wt_missionary##":"Missionär"
"##god_displeased##":"Missnöjda"
"##my_rome##":"Mitt Rom"
"##centurion_send_army_to_player##":"Mitt tålamod är slut. Då du fortfarande inte har bra relation med Kjesaren, måste jag tyvärr utföra mina order, oavsett hur otäcka de är. Ge upp nu eller bered dig på konsikvenserna!"
"##furniture_workshop##":"Möbelsnickeri"
"##furniture##":"Möbler"
"##furniture_need##":"Möbler behövs"
"##sdlr_bold##":"Modig"
"##statue_big_info##":"Monument över framstående medborgare och historiska händelser ger ett område bättre status. Folket är stolta över att ha statyer i grannskapet... och ju större desto bättre."
"##legion_morale##":"Moral"
"##native_center_info##":"Mötesplats för lokalbefolkningen"
"##nativeCenter_info##":"Mötesplatsen för den lokalbefolkning som kommer hit för att byteshandla med enkla handelsvaror. Om styresmannen bara kunde lära sig några ord på latin..."
"##wall##":"Mur"
"##walls_need_a_gatehouse##":"Murar behöver grindstugor, så att vandringsmän och handelsmän kan komma och gå som de vill."
"##fortification_info##":"Murar saktar ner fiendens framstöt mot en stad. Murar kan raseras. Tjockare murar är starkare och dessutom ges vaktposterna i anslutna torn möjlighet att patrullera dem."
"##wall_info##":"Murar skyddar värnlösa medborgare från barbarer. De kan bara motstå en viss grad av attacker, och tjockare murar klarar sig längre."
"##tooltip_some##":"Mushjälp - DELVIS"
"##tooltip_full##":"Mushjälp - FULL"
"##gmsndwnd_theme_sound##":"Musik"
"##music##":"MUSIK:"
"##god_verygood##":"Mycket bra"
"##god_quitepoor##":"Mycket dålig"
"##god_verypoor##":"Mycket dålig"
"##non_cvrg##":"Mycket dålig"
"##sld_quite_daring##":"Mycket djärv"
"##vegetable_farm_slow_work##":"Mycket få jordbrukare arbetar här. De få grönsaker som odlas är små och osunda."
"##pottery_bad_work##":"Mycket få människor arbetar här. Som resultat går krukproduktionen långsamt."
"##fig_farm_bad_work##":"Mycket få människor arbetar i denna fruktträdgård. Fruktskörden kommer att bli liten och sen."
"##weapons_workshop_slow_work##":"Mycket få människor arbetar i vapenfabriken. Som resultat är vapenproduktionen långsam."
"##meat_farm_slow_work##":"Mycket få människor arbetar på den här farmen. Som resultat är köttproduktionen långsam."
"##vinard_slow_work##":"Mycket få människor arbetar på denna odling. Som resultat är druvproduktionen långsam."
"##lumber_mill_slow_work##":"Mycket få människor arbetar vid den här brädgården. Som resultat är timmerproduktionen långsam."
"##oil_workshop_slow_work##":"Mycket få människor arbetar vid denna olivpress. Som resultat är oljeproduktionen långsam."
"##wine_workshop_slow_work##":"Mycket få människor arbetar vid denna vingård. Som resultat är vinproduktionen långsam."
"##iron_mine_slow_work##":"Mycket få människor arbetar vid det här brottet. Som resultat är järnproduktionen långsam."
"##quarry_patrly_workers##":"Mycket få människor arbetar vid det här brottet. Som resultat är marmorproduktionen långsam."
"##quarry_slow_work##":"Mycket få människor arbetar vid detta lertag. Som resultat är lerproduktionen långsam."
"##furniture_workshop_slow_work##":"Mycket få snickare arbetar här. Som resultat är möbelproduktionen långsam."
"##very_low_fire_risk##":"Mycket liten brandrisk"
"##some_defects_damage_risk##":"Mycket liten risk för kollaps"
"##sldr_very_bold##":"Mycket modig"
"##sldr_very_frightened##":"Mycket rädd"
"##very_high_fire_risk##":"Mycket stor brandrisk"
"##collapse_available_damage_risk##":"Mycket stor risk för kollaps"
"##sldr_badly_shaken##":"Mycket uppskakad"
"##middle_fest_description##":"När 1 dagsfesten närmar sig sitt slut, börjar invånare återvända hemåt, trötta men glada. Medan din valda gud ler åt dem alla."
"##military_academy_patrly_workers##":"När nya soldater har avslutat sin utbildning i förläggningen kommer de hit för att förbättra och finslipa sina färdigheter. Det går dock först när vi har fått tillräckligt med personal."
"##smcurse2_of_venus_description##":"När Venus är missnöjd sänker hon medborgarnas sinnesstämning. En del säger att hon för med sig sjukdomar."
"##wrath_of_neptune_title##":"Neptune vrede"
"##smallcurse_of_neptune_description##":"Neptunus är missnöjd med att du inte visar honom tillräcklig uppmärksamhet och frammanar en mindre storm."
"##smallcurse_of_neptune_title##":"Neptunus är upprörd"
"##smallcurse_of_neptune##":"Neptunus skyddar sjömän och deras skepp från havets faror. Om du gör honom missnöjd riskerar du dina sjömäns liv."
"##small_neptune_temple##":"Neptunustempel"
"##profit##":"Nettoflöde in/ut"
"##god_pleased##":"Nöjda"
"##north##":"Norr"
"##northBtnTooltip##":"Norr"
"##month_11_short##":"Nov"
"##lionTamer_good_life##":"Nu har du din chans, Leo. Duktigt lejon."
"##wn_numidian##":"Numidier"
"##current_play_runs_for_another##":"Nuvarande pjäs spelas i ytterligare"
"##current_game_speed_is##":"Nuvarande spelhastighet"
"##new_trade_route_to##":"Ny handelsväg etablerad."
"##plname_start_new_game##":"Ny karriär"
"##mainmenu_startcareer##":"Ny karriär"
"##mainmenu_loadmap##":"Ny karta"
"##new_map##":"Ny karta"
"##centurion_new_order_to_save_player##":"Nya order har just anlänt. Verkar som att Kjesaren har ändrat sig angående dig, och tacksamt ska jag återvända till Rom. Farväl...för denna gång."
"##newcomer_this_month##":"nykomling anlände denna månad"
"##newcomers_this_month##":"nykomlingar anlände denna månad"
"##mainmenu_newgame##":"Nytt spel"
"##ok##":"OK"
"##month_10_short##":"Okt"
"##scribemessages_unread##":"Oläst meddelande. Vänsterklicka på detta meddelande för att läsa det.  Högerklicka på detta meddelande för att radera det"
"##varieties_food_eaten##":"Olika sorters livsmedel som ätits,"
"##olive##":"Oliver"
"##olive_farm_info##":"Oliver är värdefulla för sin olja. Olivpresserierna ger olja för matlagning, belysning, smörjning och konservering."
"##olive_farm##":"Olivodling"
"##oil##":"Olja"
"##oil_workshop##":"Oljepresseri"
"##gmenu_about##":"Om"
"##romeGuard_low_entertainment##":"Om det fanns bättre underhållning i staden skulle vakttjänsten inte kännas så betungande."
"##tamer_normal_life##":"Om du rör mitt lejon, får du smaka på min piska."
"##rioter_say_3##":"Om du vill veta hur städer ser ut när de brinner, se noga på nu!"
"##warning_baths_access##":"Om ingen badhusarbetare passerar snart, kommer detta hus att förlora sin tillgång till badhus"
"##warning_barber_access##":"Om ingen barberare går förbi huset snart, kommer det att förlora sin tillgång till barberare"
"##warning_library_access##":"Om ingen bibliotekarie passerar huset snart, kommer det att förlora sin tillgång till bibliotek"
"##warning_hospital_access##":"Om ingen kirurg passerar detta hus snart, kommer det att förlora sin tillgång till sjukhus"
"##warning_doctor_access##":"Om ingen läkare passerar huset snart, kommer det att förlora sin tillgång till läkarklinik"
"##warning_college_access##":"Om ingen lärare passerar huset snart, kommer det att förlora sin tillgång till högskola"
"##warning_school_access##":"Om inget skolbarn passerar huset snart, kommer det att förlora sin tillgång till skola"
"##seamerchant_noany_trade##":"Om jag fick bestämma skulle jag inte segla den här vägen. Den här staden varken köper eller säljer något."
"##engineer_so_hungry##":"Om jag inte får mat snart ger jag mig av från staden."
"##taxCollector_gods_angry##":"Om vi inte bygger fler tempel snart, kommer gudarna att förbanna denna stad."
"##taxCollector_so_hungry##":"Om vi inte får mer livsmedel finns det snart ingen som kan betala skatt!"
"##lionTamer_so_hungry##":"Om vi inte får mer mat snart, äter lejonet upp mig!"
"##some_crime_risk##":"Området löper viss risk att drabbas av brottslighet."
"##desirability##":"Önskvärdhet"
"##open_formation_title##":"Öppen formation"
"##open_formation_text##":"Öppen ordning ger möjlighet att täcka ett brett område, men ger dem ingen formationsfördel."
"##mainmenu_randommap##":"Öppet spel "
"##fileload_load_tlp##":"Öppna detta sparade spel"
"##open_trade_route##":"Öppna handelsväg"
"##emp_open_trade_route##":"Öppna handelsväg"
"##Load_save##":"Öppna sparat spel"
"##oracle##":"Orakel"
"##oracles##":"Orakel"
"##oracles_in_city##":"Orakel i staden"
"##oracle_info##":"Orakel ökar efterfrågan på husen i stadsdelen och gör de boende gladare. Denna byggnad tillfredsställer samtliga gudar."
"##donot_organize_festival##":"Organisera ingen festival"
"##lgn_snakes##":"Ormarna"
"##east##":"Öst"
"##collapse_immitent##":"Överhängande risk för kollaps"
"##idle_factory_in_city##":"overksam industri i staden"
"##idle_factories_in_city##":"overksamma industrier i staden"
"##overlays##":"Översikt"
"##ovrm_text##":"Översikt"
"##heading_to_city_warehouses##":"På väg mot stadens handelsmagasin"
"##wt_patrician##":"Patricier"
"##egift_persian_carpets##":"Persiska mattor"
"##governor_salary_title##":"Personlig inkomst"
"##pn_salary##":"Personlig inkomst"
"##wn_picts##":"Pikter"
"##favor_rating##":"Popularitetsställning"
"##population_milestone##":"Populations milstolpe"
"##wt_priest##":"Präst"
"##miletus_win_text##":"Precis som jag förväntade mig har exemplet Miletus redan inspirerat andra östliga städer att inleda förhandlingar om att ingå i imperiet. Din erfarenhet av fisket har blivit en läxa för alla mina ståthållare!"
"##wt_prefect##":"Prefekt"
"##burning_ruins_info##":"Prefekterna kunde inte nå hit i tid för att rädda byggnaden. När elden har brunnit ut kommer endast spillror att finnas kvar på denna plats."
"##prefecture##":"Prefektur"
"##prefecture_info##":"Prefekturerna sänder prefekter till staden för att hålla fred, och för att bekämpa bränder. Ordning kan endast upprätthållas om prefekterna patrullerar staden."
"##ovrm_desirability##":"Prestige"
"##praetor_salary##":"Pretorslön på"
"##priority_level##":"Prioritetsnivå"
"##a_price_rise_title##":"Prisändringar"
"##rome_prices##":"Priser fastställs av Rom"
"##ovrm_troubles##":"Problem"
"##land_trade_problem_title##":"Problem med landhandeln"
"##rawm_production_complete_m##":"Produktionen är"
"##proconsoul_salary##":"Prokonsulslön på"
"##procurator_salary##":"Prokuratorslön på"
"##delete##":"Radera"
"##delete_this_message##":"Radera detta meddelande"
"##delete_object##":"Radera objekt"
"##delete_game##":"Radera spelet"
"##gmenu_advisors##":"Rådgivare"
"##percents##":"Ränta på"
"##god_wrathful##":"Rasande"
"##ready_to_game##":"Redo att spela"
"##advchief_religion##":"Religion"
"##ovrm_religion##":"Religion"
"##religion##":"Religion"
"##religion_in_your_city_is_flourishing##":"Religionen i din stad blomstrar. Invånarnas olika religionsbehov uppfylls, och prästerna rapporterar att gudarna är nöjda."
"##religion_advisor##":"Religiösa byggnader"
"##reservoir##":"Reservoar"
"##need_connect_to_other_reservoir##":"Reservoir bör vara ansluten till vattnetskälla"
"##ovrm_risks##":"Risker"
"##rome_need_some_goods##":"Rom är i behov av följande varor. Var snäll och skicka dem så snabbt som möjligt."
"##rome_raises_wages##":"Rom höjer lönerna"
"##rome_lowers_wages##":"Rom sänker lönerna"
"##rome_gratitude_request_text##":"Rom tackar dig för din senaste sändning. Din lojalitet skall inte glömmas."
"##try_reduce_your_salary##":"Rom tycker att din lön är för hög för din nuvarande ställning. Det skulle vara bra om du sänkte den."
"##try_reduce_your_high_salary##":"Rom tycker att din lön är för hög för din nuvarande ställning. Du borde sänka den lite."
"##barbarian_attack_text##":"Roms fiender är i utkanten av din stad. Räkna med 1 flaska vin eller 2 - och vad de mer önskar sig."
"##rotate_map_clockwise##":"Rotera kartan medurs"
"##rotate_map_counter-clockwise##":"Rotera kartan moturs"
"##rotateRightBtnTooltip##":"Rotera panel medurs"
"##rotateLeftBtnTooltip##":"Rotera panel moturs"
"##caesarea_win_text##":"Så Caesareas förre ståthållare ska alltså få behålla livet? Att rädda staden ur krisen är verkligen en bedrift. Jag kanske ska låta dig välja vilket land vi ska utvisa honom till."
"##this_year##":"Så här långt detta året"
"##year##":"Sädesmagasin lagrar"
"##years##":"Sädesmagasin lagrar"
"##lumber_mill_info##":"Såga virke för handel, eller till möbelverkstäderna. Patricierna vill ha möbler till sina villor, eller så kan du exportera det till dina handelspartners."
"##securityBtnTooltip##":"Säkerhet"
"##sell_price##":"Säljarna får"
"##emw_sold##":"Sålt"
"##citychart_society##":"Samhälle"
"##wn_samnites##":"Samniter"
"##send_modest_gift##":"Sänd en blygsam gåva"
"##send_lavish_gift##":"Sänd en frikostig gåva"
"##dispatch_gift##":"Sänd en gåva"
"##send_generous_gift##":"Sänd en generös gåva"
"##dispatch_gift_title##":"Sänd gåva till kejsaren"
"##empire_service_tip##":"Sänd iväg trupper för att skydda"
"##dispatch_force##":"Sänd iväg undsättningsstyrka?"
"##dispatch_goods?##":"Sända iväg varor?"
"##god_irriated##":"Sårade"
"##sarmizegetusa_title##":"Sarmizegetuza: en mycket farlig provins"
"##month_from_last_festival##":"sedan senaste festivalen"
"##mission_win##":"Seger"
"##sailing_to_city_docks##":"Seglar mot stadens lastkajer"
"##wn_selecids##":"Selucider"
"##senate_1##":"Senat"
"##senate##":"Senat"
"##disabled_draw_salary_for_free_reign##":"Senaten förbjuder dig att ta ut lön nu, eftersom du fortsätter att styra av egen fri vilja."
"##senate_1_info##":"Senatsbyggnaden är en av de attraktivaste byggnaderna i staden. Den ger anställning åt skatteindrivarna och inkomsterna från deras verksamhet förvaras här."
"##month_9_short##":"Sep"
"##partician_need_workers##":"Servicen blir lidande. Staden behöver fler arbetare."
"##neptune_despleasure_tip##":"Sjömän finner att Neptunus är en ombytlig gud även om han blidkas. Väck inte Neptunus vrede, om du önskar bedriva handel över vattnet."
"##hospital##":"Sjukhus"
"##hospitals##":"Sjukhus"
"##ovrm_hospital##":"Sjukhus"
"##ovrm_damage##":"Skada"
"##damage##":"Skador"
"##wt_taxCollector##":"Skatteindrivare"
"##ovrm_tax##":"Skatter"
"##tax_rate##":"Skattesatsen"
"##school##":"Skola"
"##ovrm_school##":"Skola"
"##scholar##":"Skolbarn"
"##schools##":"Skolor"
"##hlth_care_of##":"Sköter om"
"##gmspdwnd_scroll_speed##":"Skrollningshastighet"
"##stop_warehouse_devastation##":"SLUTA tömma magasin"
"##stop_granary_devastation##":"Sluta tömma sädesmagasin"
"##small_temples##":"Små tempel"
"##bldm_temple##":"Små tempel"
"##furniture_workshop_info##":"Snickarna vid snickeriet skapar fina möbler av virke. Medborgarna kan möblera sina villor och du kan handla med överskottet."
"##soldier##":"Soldat"
"##soldiers##":"Soldater"
"##soldiers_in_legion##":"Soldater i legion"
"##soldiers_health##":"Soldaternas hälsa"
"##savedlg_continue##":"Spara"
"##gmspdwnd_autosave_interval##":"Spara automatiskt"
"##save_game_here##":"Spara det aktuella spelet till denna fil"
"##dn##":"Spara karta"
"##save_map##":"Spara karta"
"##gmenu_file_save##":"Spara spel"
"##save_city##":"Spara spel"
"##special_orders##":"Specialorder"
"##game_is_paused##":"Spelet pausat (Tryck P för att fortsätta)"
"##gmspdwnd_game_speed##":"Spelhastighet"
"##operations_manager##":"Spelproducent"
"##spear##":"Spjut"
"##wt_romeSpearman##":"Spjutkastare"
"##mainmenu_language##":"Språk"
"##crack##":"Spricka"
"##rift_info##":"Sprickor i marken"
"##delivery_boy##":"Springpojke"
"##city_still_in_debt##":"Stad fortfarande i skuld"
"##city_in_debt##":"Stad i skuld"
"##city_in_debt_again##":"Stad i skuld igen"
"##cartPusher_good_life##":"Stad som stad... Den här verkar rätt bra."
"##city_options##":"Stadalternativ"
"##city_is_besieged##":"Staden är belägrad"
"##doctor_low_entertainment##":"Staden är så trist att mina patienter frågar om jag kan bota kronisk uttråkning!"
"##advchief_workless##":"Staden har en arbetslöshet på"
"##advchief_employers_ok##":"Staden har inga arbetslöshetsproblem"
"##advchief_needworkers##":"Staden saknar"
"##taxCollector_average_life##":"Staden tycks fungera väl."
"##city_have_defence##":"Stadens försvar skulle aldrig ha släppt igenom fienden!"
"##advchief_health_high##":"Stadens hälsosituation är bra"
"##advchief_health_high_clinic##":"Stadens hälsosituation är bra, dina medborgare lider bara av enklare sjukdomar."
"##advchief_health_bad##":"Stadens hälsosituation är dålig"
"##advchief_health_bad_clinic##":"Stadens hälsosituation är dålig, dina överansträngda läkare fruktar en dödlig epidemi."
"##advchief_health_less_clinic##":"Stadens hälsosituation är dålig, mat och kliniker skulle förbättra hälsan."
"##advchief_health_low##":"Stadens hälsosituation är förfärande"
"##advchief_health_lower##":"Stadens hälsosituation är förfärande, pest kommer med all säkerhet bryta ut."
"##advchief_health_terrible##":"Stadens hälsosituation är fruktansvärd"
"##advchief_health_terrible_clinic##":"Stadens hälsosituation är fruktansvärd, klinikerna hinner inte med, sjukdomar är nästan oundvikliga."
"##advchief_health_less##":"Stadens hälsosituation är ganska dålig"
"##advchief_health_simple##":"Stadens hälsosituation är inte bra, se till att dina medborgare har mat och kliniker."
"##advchief_health_simple_clinic##":"Stadens hälsosituation är mindre bra"
"##advchief_health_verygood##":"Stadens hälsosituation är mycket bra"
"##advchief_health_verygood_clinic##":"Stadens hälsosituation är mycket bra, medborgarnas småkrämpor hanteras snabbt av lokala läkare."
"##advchief_health_good##":"Stadens hälsosituation är nästan perfekt"
"##advchief_health_good_clinic##":"Stadens hälsosituation är nästan perfekt, läkarnas kliniker är nästan tomma."
"##advchief_health_perfect##":"Stadens hälsosituation är perfekt"
"##advchief_health_perfect_clinic##":"Stadens hälsosituation är perfekt, dina tomma kliniker utgör ett exempel genom hela imperiet."
"##advchief_health_middle##":"Stadens hälsosituation är tillfredsställande"
"##advchief_health_middle_clinic##":"Stadens hälsosituation är tillfredsställande, klinikerna håller farliga epidemier borta."
"##advchief_health_awesome_clinic##":"Stadens hälsosituation är utmärkt, inga väntetider alls för besök till lokala läkare."
"##advchief_health_awesome##":"Stadens hälsosituation är utmärkt."
"##doctor_good_life##":"Stadens invånare tycks vara vid god hälsa."
"##city_settings##":"Stadinställningar"
"##rating##":"Ställning"
"##wnd_ratings_title##":"Ställning"
"##how_to_grow_prosperity##":"Ställningen har inte förändrats detta året. Att visa vinst i stadens årliga räkenskaper är det bästa sättet att förbättra välståndsställningen."
"##advchief_sentiment##":"Stämning"
"##poor_city_mood_lack_migration##":"Stämningen i staden förhindrar immigration"
"##close##":"Stäng"
"##infobox_tooltip_exit##":"Stäng detta fönster"
"##sldh_health_strong##":"Stark"
"##tradeadv_industrystate_tip##":"Starta eller avsluta produktion för denna aktivitet överallt i staden"
"##gmenu_file_restart##":"Starta om"
"##need_restart_for_apply_changes##":"Starta om spelet för att aktivera de nya inställningarna"
"##start_condition##":"Startvillkor"
"##rioter_say_1##":"Ståthållaren bryr sig uppenbarligen inte om mig, så jag tänker visa vad jag tycker om hans stad."
"##valentia_preview_mission##":"Ståthållaren ställs inför olika hot och faror, och Iberierna utgör inte det minsta av dessa! De har inte för avsikt att ge upp Hispanien."
"##governor_palace_1##":"Ståthållarens hus"
"##governorHouse##":"Ståthållarens hus"
"##governor_palace_3##":"Ståthållarens palats"
"##governorPalace##":"Ståthållarens palats"
"##governor_palace_2##":"Ståthållarens villa"
"##governorVilla##":"Ståthållarens villa"
"##fort_horse##":"Stödtrupp - Ridande"
"##high_fire_risk##":"Stor brandrisk"
"##middle_festival##":"Stor festival"
"##big_shack##":"Stor koja"
"##advchief_high_crime##":"Stor kriminalitet råder i staden"
"##high_damage_risk##":"Stor risk att kollapsa"
"##statue_big##":"Stor staty"
"##beatifull_villa##":"Stor villa"
"##large_temples##":"Stora tempel"
"##bldm_big_temple##":"Stora tempel"
"##great_festival##":"Storslagen festival"
"##beatyfull_insula##":"Storslagen Insulae"
"##large##":"Stort"
"##big_hovel##":"Stort skjul"
"##large_temple##":"Stort tempel"
"##difficulty##":"Svårighetsgrad"
"##lgn_pigs##":"Svinen"
"##meat_farm##":"Svinuppfödning"
"##south##":"Syd"
"##southEast##":"Sydost"
"##southWest##":"Sydväst"
"##syracusae_title##":"Syracusae: en något farlig provins"
"##destroy_bridge_warning##":"Ta ned broar med försiktighet. Isolerade samhällen kommer försvinna utan tillgång till huvudvägen till Rom."
"##thanks_to##":"TACK TILL:"
"##carthago_win_text##":"Tack vare din briljanta insats ligger det karthagiska hotet äntligen bakom oss. Våra forna fiender är nu laglydiga romerska medborgare. I alla fall de som ännu är i livet!"
"##coverage##":"Täckning i staden"
"##house_provide_food_themselves##":"Tältboende hämtar sin egen mat från omgivande marker."
"##tarentum_title##":"Tarente: une petite province dangereuse"
"##tarentum_slightly_dangerous_province##":"Tarentum: en inte helt ofarlig provins"
"##tarraco_title##":"Tarraco: en fredlig provins"
"##tarraco_win_text##":"Tarracos livsmedelsexport hjälpte imperiet att överleva en svår period. Medborgarna är skyldiga dig för sina liv och ståthållarna sina arbeten. Skördarna blir nu normala igen och jag vill använda dina talanger inom ett nytt område."
"##tarsus_title##":"Tarsus: en mestadels fredlig provins"
"##house_pay_tax##":"Taxbetalande hus"
"##theater##":"Teater"
"##ovrm_theater##":"Teatrar"
"##theaters##":"Teatrar"
"##theater_need_actors##":"Teatrarna och amfiteatrarna söker alltid efter nya talanger."
"##mainmenu_dlc_soundtrack##":"Teman"
"##temples##":"Tempel"
"##templeBtnTooltip##":"Tempel"
"##testers##":"TESTARE:"
"##time_since_last_gift##":"Tid sedan senaste gåva"
"##to_trade_advisor##":"Till handelsrådgivaren"
"##to_empire_road##":"Till Imperiet"
"##to_rome_road##":"Till Rom"
"##mission_wnd_tocity##":"Till staden"
"##dedicate_fectival_ceres##":"Tillägna Ceres en festival"
"##dedicate_fectival_mars##":"Tillägna Mars en festival"
"##dedicate_fectival_mercury##":"Tillägna Merkurius en festival"
"##dedicate_fectival_neptune##":"Tillägna Neptunus en festival"
"##dedicate_fectival_venus##":"Tillägna Venus en festival"
"##have_no_access_to_library##":"Tillgång till bibliotek krävs nu i vissa delar av staden. Dina medborgare har tid att läsa. Nu behöver de tillgång till litteratur."
"##timber##":"Timmer"
"##tingis_title##":"Tingis: en farlig provins"
"##infobox_construction_comma_tip##":"TIPS: Använd komma och punkt för snabbflyttning genom dessa och andra objekt."
"##missionBtnTooltip##":"Titel på provinskarta."
"##devastate_granary##":"Töm sädesmagasin"
"##plaza_caption##":"Torg"
"##plaza##":"Torg"
"##trees_and_forest_caption##":"Träd och skogsland"
"##trees_and_forest_text##":"Träden kan inte forceras, men de kan röjas undan. De är livsviktiga för skogsindustrin, brädgårdar måste ligga nära träden för att producera timmer."
"##garden##":"Trädgårdar"
"##gardens_info##":"Trädgårdar förbättrar den lokala miljön."
"##empire_tax##":"Tribut"
"##triumphal_arch##":"Triumfbåge"
"##wrath_of_venus_description##":"Tyvärr för dina olyckliga medborgare, Venus har inget annat val än att dela sin olycka, sprider sjukdom och elände hela folket."
"##warehouse_low_personal_warning##":"Underbemannad. Kan endast sända iväg varor, ej ta emot varor"
"##max_available##":"Underhåller"
"##entertainment_short##":"Underhållning"
"##advchief_entertainment##":"Underhållning"
"##entertainment##":"Underhållning"
"##ovrm_entertainments##":"Underhållning"
"##entertainmentBtnTooltip##":"Underhållning"
"##new_ruler##":"Une nouvelle règle"
"##showing_agamemnon_aeschylus##":"Uppför: 'Annales', av Tacitus"
"##showing_thecrito_plato##":"Uppför: 'Oidipus', av Sofokles"
"##showing_odyssey_homer##":"Uppför: 'Platons filosofi'"
"##showing_lisistrata_aristopanes##":"Uppför: 'Vergilius dikter'"
"##showing_antigone_sophocles##":"Uppför: Homeros grekiska tragedier"
"##last_riots_bad_for_peace_rating##":"Upploppen som nyligen ägde rum i staden har haft negativ inverkan på din fredsställning!"
"##fullscreen_off##":"Upplösning"
"##sldr_encouraged##":"Uppmuntrad"
"##mopup_formation_title##":"Upprensningsformation"
"##wt_rioter##":"Upprorsman"
"##sldr_shaken##":"Uppskakad"
"##original_game##":"URSPRUNGLIGA SPELET:"
"##tower_no_workers##":"Utan bemanning har vi ingen personal till våra katapulter eller vakter som kan patrullera murarna."
"##forum_no_workers##":"Utan indrivare bidrar det här kontoret inte med någonting till stadskassan."
"##prefecture_no_workers##":"Utan personal blir den här stationen inte mycket mer än en måltavla för vandaler."
"##lion_pit_no_workers##":"Utan personal kan detta lejonhus inte leverera några nya lejon till spelen."
"##gladiator_pit_no_workers##":"Utan utbildningspersonal kan denna skola inte utbilda nya gladiatorer."
"##advchief_education##":"Utbildning"
"##education_advisor_title##":"Utbildning"
"##education##":"Utbildning"
"##educationBtnTooltip##":"Utbildning"
"##ovrm_educations##":"Utbildning"
"##education_objects##":"Utbildningsbyggnader"
"##credit##":"Utgifter"
"##god_excellent##":"Utmärkt"
"##freespace_for##":"Utrymme för"
"##exit_point##":"Utträdespunkt"
"##developers##":"UTVECKLARE:"
"##healthadv_some_regions_need_hospital##":"Utvecklingen i vissa områden hålls tillbaka av för få sjukhus i staden. Nya sjukhus attraherar fler patricierklasser till staden."
"##road_caption##":"Väg"
"##road_text##":"Vägarna är livsviktiga för stadens funktion. Invånarna går bara ut ur sina hus om det finns en väg."
"##wt_cartPusher##":"Vagndragare"
"##roadBlock##":"Vägstopp"
"##wt_romeGuard##":"Vaktpost"
"##valencia_title##":"Valentia: en relativt fredlig provins"
"##select_location##":"Välj destination"
"##select_this_graph##":"Välj detta diagram"
"##select_city_layer##":"Välj en översiktsrapport för staden"
"##enter_your_name##":"Välj ett namn"
"##meat_farm_info##":"Välmående medborgare njuter av olika sorters fläsk. Kött kan förvaras i sädesmagasin för lokal konsumtion eller i handelsmagasin för export."
"##senatepp_prsp_rating##":"Välstånd"
"##wndrt_prosperity##":"Välstånd"
"##rioter_in_city_text##":"Vandalism i staden"
"##rioter_in_city_title##":"Vandalism i staden"
"##left_click_open_right_erase##":"Vänsterklicka på ett meddelande för att läsa. Högerklicka för att radera."
"##weapon##":"Vapen"
"##weapons_workshop_info##":"Vapensmeder förvandlar järn till vapen och rustningar, som du kan handla med och göra vinst eller använda för att utrusta dina egna legioner."
"##weapons_workshop##":"Vapensmedja"
"##weapon_store_of##":"Vapenupplaget har"
"##wharf_our_boat_return##":"Vår båt seglar mot hamn."
"##wharf_our_boat_fishing##":"Vår fiskebåt befinner sig vid fiskevattnet och fångar just nu fisk."
"##no_fishplace_in_city##":"Vår fiskebåt hoppas snart kunna hitta en fiskeplats. Det blir svårt att försörja sig om vi inte hittar fisk..."
"##wharf_out_boat_return_with_fish##":"Vår fiskebåt seglar tillbaka från fiskevattnen med sin fångst."
"##wharf_out_boat_ready_fishing##":"Vår fiskebåt seglar ut till fiskevattnen."
"##gladiator_gods_angry##":"Var hälsad, medborgare. Har du hört? Gudarna är vreda."
"##engineer_good_life##":"Var hälsad! Är det inte en fantastisk stad?"
"##taxCollector_good_life##":"Var hälsad! Detta är en mycket trevlig stad att bo i."
"##recruter_high_workless##":"Var hälsad! Har du sett hur hög arbetslösheten är?"
"##marketKid_say_3##":"Var hälsad! Jag bär korgen med mat till kvinnans marknad. Jag hoppas jag får bra med dricks!"
"##wt_missioner_average_life##":"Var hälsad! Jag ser att det finns mycket att göra med att lära dessa barbarer fördelarna med Roms välvilja."
"##recruter_good_life##":"Var hälsad! Livet här är gott."
"##missioner_high_barbarian_risk##":"Var hälsad! Min undervisning om Roms välvilja tycks tränga in hos dessa ganska skrämmande barbarer."
"##lionTamer_good_education##":"Var hälsad. Den här staden tycker vi om, inte sant, Leo?"
"##priest_so_hungry##":"Var hälsad. Denna stad behöver omedelbart mer livsmedel."
"##recruter_normal_life##":"Var hälsad. Detta är en ganska bra stad."
"##gladiator_good_life##":"Var hälsad. Livet här är skönt att leva, inte sant?"
"##partician_good_life##":"Var hälsad. Staden sköts riktigt bra."
"##forum_1_on_patrol##":"Vår indrivare är ute på inspektion."
"##forum_1_ready_for_work##":"Vår indrivare förbereder sig för att ge sig av."
"##engineering_post_on_patrol##":"Vår ingenjör är ute och arbetar."
"##engineering_post_ready_for_work##":"Vår ingenjör förbereder sig för att ge sig av."
"##out_legion_go_to_location##":"Vår legion marscherar för att rädda en av rikets städer"
"##out_legion_back_to_city##":"Vår legion marscherar tillbaka till vår stad"
"##prefecture_on_patrol##":"Vår prefekt är ute och patrullerar."
"##prefecture_ready_for_work##":"Vår prefekt förbereder sig för sin tjänst."
"##empiremap_our_city##":"Vår stad!"
"##dock_cart_wait##":"Vår vagn är här och väntar på nya order."
"##dock_cart_taking_goods##":"Vår vagn för varorna till annan plats."
"##our_enemies_near_city##":"Våra fiender är inom synhåll från staden"
"##our_foods_level_are_low##":"Våra livsmedelsförråd är små"
"##market_about##":"Våra marknader gör imperiets rika håvor tillgängliga för medborgare med pengar. Varje hem behöver tillgång till en marknad, men ingen vill bo intill en."
"##wt_wolf##":"Varg"
"##lgn_wolves##":"Vargarna"
"##warehouse_full_warning##":"VARNING Denna lagerbyggnad är helt fylld. Den kan inte ta emot fler varor."
"##warehouse_gettinfull_warning##":"VARNING Denna lagerbyggnad håller på att bli full. Den kan bara ta emot varor som redan finns, inga nya varutyper."
"##changesalary_greater_salary##":"Varning: Betala dig själv en lön som överstiger din grad imponerar inte på kejsaren."
"##working_build_poor_labor_warning##":"Varning: Dålig tillgång till arbetskraft"
"##working_building_need_road##":"VARNING. Denna byggnad fungerar ej. Den ligger inte intill en väg, och dess anställda kommer ej fram"
"##warning_some##":"Varningar AV"
"##warning_full##":"Varningar PÅ"
"##city_warnings_off##":"Varningar: Av"
"##city_warnings_on##":"Varningar: På"
"##warehouse_info##":"Varor som produceras för handel kräver magasinering. Karavaner besöker handelsmagasinen för att köpa och sälja varor och handelshamnar får sitt gods från intilliggande magasin."
"##cartPusher_need_workers##":"Vart man än kommer i staden finns det lediga arbeten."
"##west##":"Väst"
"##ovrm_water##":"Vatten"
"##water_caption##":"Vatten"
"##water_supply##":"Vatten"
"##show_spots_of_city_troubles_tip##":"Växla mellan aktuella problemområden i staden"
"##venus##":"Venus"
"##smcurse_of_venus_title##":"Venus är upprörd"
"##blessing_of_venus_description##":"Venus förmedlar en känsla av välvilja till din stad, vilket får alla dina medborgare på bättre humör."
"##wrath_of_venus_title##":"Venus vrede"
"##smcurse_of_venus_description##":"Venus, förmedlare av kärlek och harmoni, är upprörd. Detta bådar inget gott för prefekterna i din stad!"
"##small_venus_temple##":"Venustempel"
"##emigrant_high_workless##":"Vet ni var det kan finnas arbete? Jag måste få ett arbete."
"##wheat##":"Vete"
"##wheat_farm_info##":"Vetekorn är det grundläggande livsmedlet för ditt folk. Det måste lagras i sädesmagasin för att livnära ditt folk, eller i handelsmagasin för export."
"##wheat_farm##":"Veteodling"
"##sldr_totally_distraught##":"Vettskrämd"
"##forum_1_slow_work##":"Vi är kraftigt underbemannade och har en lucka på två veckor innan indrivarna ger sig ut."
"##engineering_post_slow_work##":"Vi är kraftigt underbemannade och har en tidslucka på två veckor mellan ingenjörernas rundor."
"##lion_pit_need_some_workers##":"Vi är något underbemannade, och kan därför endast leverera två nya lejon i månaden."
"##gladiator_pit_need_some_workers##":"Vi är något underbemannade, och kan därför endast utbilda två nya gladiatorer i månaden."
"##dock_need_some_workers##":"Vi är underbemannade och därför kommer det att ta lite längre tid än vanligt att lasta och lossa de fartyg som anlöper hamnen."
"##forum_patrly_workers##":"Vi är underbemannade och måste vänta en vecka innan våra indrivare är tillbaka i tjänst."
"##barracks_bad_weapons_slow_workers##":"Vi är underbemannade och saknar vapen, vi kan bara långsamt utbilda stödtrupper."
"##barracks_have_weapons_slow_workers##":"Vi är underbemannade och utbildar nya soldater långsamt, men vi har de vapen som krävs för att utbilda alla typer av soldater."
"##prefecture_patrly_workers##":"Vi är underbemannade, och har farliga luckor på upp till en vecka i vår tjänstgöringslista."
"##prefecture_bad_work##":"Vi arbetar endast med kontorspersonal. Det går ofta en hel månad utan att vi sänder en prefekt ut på gatorna."
"##engineering_post_bad_work##":"Vi arbetar med minimistyrka. Vi kan knappt sända ut en ingenjör per månad på fältet."
"##missionaryPost_full_work##":"Vi arbetar på att civilisera lokalbefolkningen. Genom att lära dem grunderna i latin hoppas vi uppmuntra dem att arbeta med oss, istället för emot oss."
"##we_eat_more_thie_produce##":"Vi äter mer än vi producerar"
"##we_eat_much_then_produce##":"Vi äter mycket mer än vi producerar"
"##we_eat_some_then_produce##":"Vi äter något mer än vi producerar"
"##dock_busy_bad_work##":"Vi betjänar det förtöjda fartyget, men har för få hamnarbetare, detta kommer att ta tid."
"##dock_busy_patrly_workers##":"Vi betjänar det förtöjda fartyget, trots att vi inte har tillräckligt med anställda, så det kommer att ta längre tid än det borde."
"##getting_reports_about_enemies##":"Vi får rapporter om fiender som närmar sig staden"
"##restocking_fishing_boat##":"Vi förbereder för närvarande vår fiskebåt för att segla ut igen. Hur snabbt det går beror på hur många anställda vi har."
"##militaryAcademy_full_work##":"Vi förser nya rekryter från stadens förläggningar med den ytterligare utbildning de kräver för att fungera bra i en modern romersk armé."
"##prefecture_slow_work##":"Vi har alldeles för få prefekter. Det händer att inga prefekter lämnar stationen på upp till två veckor åt gången."
"##lion_pit_patrly_workers##":"Vi har bara halva personalstyrkan, och kan därför endast leverera ett lejon under nästa månad."
"##gladiator_pit_patrly_workers##":"Vi har bara halva personalstyrkan, och kan därför endast utbilda en gladiator under nästa månad."
"##engineering_post_patrly_workers##":"Vi har för lite personal, så vi måste vänta en vecka innan våra ingenjörer är tillbaka i tjänst."
"##dock_full_work##":"Vi har full arbetsstyrka och kommer att kunna lasta och lossa inkommande fartyg."
"##dock_no_workers##":"Vi har inga hamnarbetare och kan därför inte lasta eller lossa några fartyg som kommer till hamnen."
"##no_warning_for_us##":"Vi har inga rapporter om hot"
"##forum_need_some_workers##":"Vi har korta avbrott i verksamheten, ungefär en dag eller två, innan våra indrivare är tillbaka på gatorna igen."
"##prefecture_need_some_workers##":"Vi har lite ont om prefekter. Vi har luckor på en dag eller två i vår täckning."
"##dock_bad_work##":"Vi har mycket få hamnarbetare så det kommer att ta lång tid att lasta och lossa de fartyg som anlöper hamnen."
"##tower_have_workers_no_soldiers##":"Vi har underhållspersonal, men vi behöver trupper från en förläggning för att försvara staden."
"##barracks_no_weapons##":"Vi kan utbilda stödtrupper mycket snabbt, men utan vapenupplag kan vi inte utbilda några nya legionärer."
"##lion_pit_slow_work##":"Vi lider av svår personalbrist, och kommer att få kämpa för att leverera ett enda lejon under de kommande två månaderna."
"##gladiator_pit_slow_work##":"Vi lider av svår personalbrist, och kommer att få kämpa för att utbilda en ny gladiator under de kommande två månaderna."
"##we_produce_some_than_eat##":"Vi producerar lagom för att livnära alla"
"##we_produce_much_than_eat##":"Vi producerar mycket mer än vi äter"
"##we_produce_more_than_eat##":"Vi producerar något mer än vi äter"
"##barracks_bad_weapons_need_some_workers##":"Vi saknar några anställda och utbildar soldater långsammare än vanligt. Utan vapenupplag kan vi inte utbilda några nya legionärer."
"##enemies_very_hard##":"Vi ska göra vårt bästa, men även romerska soldater får svårt att besegra den här fienden."
"##enemies_very_easy##":"Vi ska nog skrämma bort veklingarna snabbt."
"##barracks_city_not_need_soldiers##":"Vi utbildar för närvarande inga rekryter eftersom vi inte har fått någon begäran från stadens fort eller torn om nya styrkor."
"##wait_for_fishing_boat##":"Vi vänta för närvarande på att ett varv skall bygga oss en fiskebåt."
"##londinium_win_text##":"Vid Jupiter! Vildarna i Britannia har aldrig sett Londiniums like. Claudius, som visade öborna de romerska svärdens vassa eggar för många år sedan, ler säkert mot oss från sin himmel."
"##wine##":"Vin"
"##theater_no_workers##":"Vinden är det enda som rör sig i denna teater. Utan arbetare erbjuder den inga pjäser till lokalbefolkningen."
"##grape##":"Vindruvor"
"##wine_workshop##":"Vingård"
"##wine_workshop_info##":"Vinhandlare förvandlar druvor till vin, vilket patricierna kräver om de skall bygga villor. Vin är en handelsvara som är begärlig för många."
"##winning_population##":"Vinnande befolkning"
"##maximizeBtnTooltip##":"Visa fönster"
"##show_bigpanel##":"Visa hela sidopanelen"
"##infobox_tooltip_help##":"Visa hjälpen för detta fönster"
"##show_prices##":"Visa priser"
"##wn_visigoth##":"Visigoter"
"##some_fire_risk##":"Viss brandrisk"
"##little_damage_risk##":"Viss risk att kollapsa"
"##some_amphitheaters_no_actors##":"Vissa av dina amfiteatrar saknar skådespelare och gladiatorer. Fler underhållare skulle ge bättre villkor i de stadsdelar som klagar över dålig underhållning."
"##healthadv_some_regions_need_doctors##":"Vissa delar av staden kräver tillgång till en klinik. Utan någon form av hälsovård kommer dessa hus förmodligen inte att växa."
"##healthadv_some_regions_need_bath##":"Vissa delar av staden vill ha fler badhus. Vissa hus har tillgång till bad, men andra har det inte, och detta hindrar deras utveckling."
"##advchief_some_need_baths##":"Vissa medborgare behöver badhus"
"##advchief_some_need_barber##":"Vissa medborgare behöver barberare"
"##advchief_some_need_doctors##":"Vissa medborgare behöver läkarkliniker"
"##advchief_some_need_hospital##":"Vissa medborgare behöver sjukhus"
"##some_houses_need_amph_for_grow##":"Vissa medborgare klagar över bristande tillgång till fritidsanläggningar. Vissa områden i staden kräver mer varierade underhållningsmöjligheter."
"##some_houses_inadequate_entertainment##":"Vissa medborgare klagar över bristande tillgång till underhållning i sina områden. Du kanske behöver erbjuda ett mer varierat utbud, eller kanske bygga fler skådespelarkolonier till dina teatrar."
"##religionadv_need_third_religion##":"Vissa medborgare vill ha en tredje religion etablerad nära sitt område. De anser att detta skulle attrahera bättre patricierklasser."
"##advchief_some_need_library##":"Vissa medborgare vill ha fler bibliotek"
"##advchief_some_need_academy##":"Vissa medborgare vill ha fler skolor"
"##advchief_high_crime_in_district##":"Vissa områden har hög kriminalitet"
"##advchief_which_crime_in_district##":"Vissa områden har mindre problem"
"##healthadv_some_regions_need_bath_2##":"Vissa områden i staden behöver nu tillgång till badhus. Bristen på dessa sanitära anläggningar begränsar byggnadstillväxten i dessa områden."
"##some_houses_need_library_or_colege_access##":"Vissa områden i staden kräver nu skolor och högskolor. Bristen på utbildningsmöjligheter förhindrar byggandet av bättre bostäder i dessa områden."
"##some_houses_need_better_library_access##":"Vissa områden i staden vill ha bättre tillgång till bibliotek. Välbärgade medborgare tycker om att läsa men vill inte gå långt för att nå biblioteket."
"##have_no_access_school_colege##":"Vissa områden kräver bättre tillgång till skolor och högskolor. Endast vissa hus har tillgång till skolor eller högskolor, och detta hindrar områdenas utveckling."
"##nativeField_info##":"Vissa primitiva grödor, som förser lokalbefolkningen med en grundläggande källa till livsmedel."
"##some_soldiers_need_weapon##":"Vissa soldater måste ha tillgång till vapenförråd"
"##healthadv_some_regions_need_barbers_2##":"Vissa välbeställda delar av staden vill ha barberare. En lokal barberare ger bättre status åt området."
"##gmsndwnd_game_volume##":"Volym"
"##floatsam##":"Vrakgods"
"##floatsam_enabled##":"Vrakgods på?"
"##god_veryangry##":"Vredgade"
"##city_zoom_off##":"Zoom: Av"
"##city_zoom_on##":"Zoom: På"
"##procurator##":"Procurator"
"##proconsul##":"Proconsul"
"##praetor##":"Praetor"
"##spirit_of_mars_text##":"Andan väktare trollade av Mars för att skydda dig vaknar, och lägger låg några av dem som vågar angripa hans valda staden."
"##smallcurse_of_mars_failed_text##":"Mars är vrede med dig. Skratta om du inte är rädd, eftersom även idag kan du inte föra krig, kommer Mars inte glömma förolämpningar tillfogat honom. Akta dig!"
}