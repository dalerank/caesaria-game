{"##some_food_on_next_month##":"- vissa livsmedel till kommande månad",
"##have_no_food_on_next_month##":"- inga livsmedel till kommande månad",
"##small_food_on_next_month##":"- mycket lite mat till kommande månad",
"##city_barbarian_off_tlp##":"Barbarer kommer inte attakera din stad",
"##city_barbarian_off##":"Barbarer: AV",
"##city_barbarian_on##":"Barbarer: ON",
"##city_barbarian_on_tlp##":"Barbarer kan komma attackera din stad",
"##city_c3rules_off_tlp##":"Spelet använder reglerna från Caesar III och nya",
"##city_c3rules_off##":"C3 regler + nya regler",
"##city_c3rules_on##":"C3 regler bara",
"##city_df_usual_tlp##":"Normal svårighetsgrad, brott och skatter",
"##city_df_hard_tlp##":"Ökadade risker för upplopp, lägre skatter
",
"##city_df_fun_tlp##":"Inga upplopp i staden, mindre påverkan av gudar, skatter opåverkade",
"##city_df_easy_tlp##":"Liten risk för uppror, höga skatter, nästan ingen påverkan från gudarna",
"##city_df_simple_tlp##":"Normal risk för uppror, ingen korruption, normala skatter",
"##city_df_usual##":"Normal svårighetsgrad",
"##city_df_hard##":"Ökad svårighetsgrad
",
"##city_df_nicety##":"Mycket hög svårighetsgrad",
"##city_df_impossible##":"Omöjligt",
"##city_df_fun##":"För skoj skull",
"##city_df_easy##":"Lätt svårighetsgrad",
"##city_df_simple##":"Enkelt att spela",
"##city_opts_god_on_tlp##":"Gudarna påverkar livet i staden",
"##city_opts_god_off_tlp##":"Gudarna är inte intresserade av din stad",
"##city_chastener_on_tlp##":"Caesar kan skicka dödspatrullen",
"##city_chastener_off_tlp##":"Caesar kommer inte skicka dödspatrullen",
"##city_chastener_on##":"Caesar legion: PÅ",
"##city_chastener_off##":"Caesar legion: AV",
"##city_androidbar_on_tlp##":"Visa fönstret för mobilenheter",
"##city_androidbar_off_tlp##":"Fönstret för mobilaenheter visas inte",
"##city_androidbar_on##":"Adv. alternativ: VISA",
"##city_androidbar_off##":"Adv. alternativ: Dölj",
"##city_debug_on_tlp##":"Debugmeny tillgänglig",
"##city_debug_off_tlp##":"Debugmeny dold",
"##city_debug_on##":"Debugmeny: VISA",
"##city_debug_off##":"Debugmeny: DÖLJ",
"##city_destroy_epdh_off_tlp##":"Staden påverkas inte av epedimier",
"##city_destroy_epdh_on_tlp##":"Staden påverkas av epedimier",
"##city_forest_fire_on_tlp##":"Skogen kan fatta eld
",
"##city_forest_fire_off_tlp##":"Skogen kan inte fatta eld
",
"##city_forest_grow_off_tlp##":"Skogen vill inte växa",
"##city_forest_grow_on_tlp##":"Skogen kan växa",
"##city_destroy_epdh_off##":"Ext. epidemi regler",
"##city_destroy_epdh_on##":"Enkla epidemi regler
",
"##city_forest_fire_on##":"Skogsbränder: På",
"##city_forest_fire_off##":"Skogsbränder: Av",
"##city_forest_grow_off##":"Skogen växer: Av",
"##city_forest_grow_on##":"Skogen växer: På",
"##city_zoominv_on_tlp##":"Normalzoom",
"##city_zoominv_off_tlp##":"Inveterad normalzoom",
"##city_lockinfo_on_tlp##":"Infofönster kan inte flyttas",
"##city_lockinfo_off_tlp##":"Infofönster kan flyttas",
"##city_mapmoving_lmb_tlp##":"Flytta runt kartan genom att hålla ned vänster musknapp",
"##city_mapmoving_mmb_tlp##":"Flytta runt kartan genom att hålla ned mittersta musknappen",
"##city_tooltips_on_tlp##":"Visa tips i staden",
"##city_tooltips_off_tlp##":"Visa inte tips i staden",
"##city_lockinfo_on##":"Infofönster: LÅST",
"##city_lockinfo_off##":"Infofönster: FLYTTAD",
"##city_mapmoving_lmb##":"Flytta kartan: vänster musknapp",
"##city_mapmoving_mmb##":"Flytta kartan: mittersta musknappen",
"##city_tooltips_on##":"Visa tips: PÅ",
"##city_tooltips_off##":"Visa tips: AV",
"##city_warnings_on_tlp##":"Inkludera debugmeddelanden",
"##city_warnings_off_tlp##":"Inkludera inte debugmeddelanden",
"##city_zoom_on_tlp##":"Zoom är aktivt",
"##city_zoom_off_tlp##":"Zoom inte aktivt",
"##dn_for_open_trade##":"för att öppna handelsväg",
"##target_population_is##":"( Målbefolkningen är",
"##no_target_population##":"( Ingen målbefolkning )",
"##mainmenu_mcmxcviii##":"MCMXCVIII",
"Variable":"SVENSKA (v1.0)",
"##age_uc##":"UC",
"##actor_gods_angry##":"Aaagh!! Gudarna är rasande. Vi går under!",
"##ovrm_aborigen##":"Aborigin",
"##month_8_short##":"Ago",
"##mainmenu_credits##":"Credits",
"##extm_administration_tlp##":"Administrativa- eller regeringsbyggnader",
"##ovrm_academy##":"Högskola",
"##colleges##":"Högskolor",
"##academy##":"Högskola",
"##aqueduct##":"Akvedukt",
"##aqueduct_info##":"Akvedukter gör det möjligt att konstruera reservoarer långt från vatten, vilket gör det möjligt för fontäner att förse staden med vatten.",
"##actor##":"Skådespelare",
"##advchief_haveprofit##
":"Tillgångarna har i år stigit med",
"##advchief_havedeficit##":"Tillgångarna har i år minskat med",
"##granery##":"Sädesmagasin",
"##granary_holds##":"Sädesmagasin innehåller
",
"##granaries_holds##":"Sädesmagasiner innehåller
",
"##amphitheater##":"Amfiteater",
"##amphitheatres##":"Amfiteatrar",
"##ovrm_amphitheater##":"Amfiteatrar",
"##amphitheaters##":"Amfiteatrar",
"##month_4_short##":"Apr",
"##arabian_stallions##":"Arabiska hingstar",
"##architect##":"Arkitekt",
"##balance##":"Balans",
"##ballista##":"Katapult",
"##ovrm_baths##":"Bad",
"##baths##":"Badhus",
"##bathlady##":"Badarbetare",
"##bath_1##":"Badhus",
"##bath##":"Badhus",
"##tower_may_build_on_thick_walls##":"Du kan endast bygga torn på tjocka murar",
"##tower##":"Torn",
"##engineering_post_no_workers##":"Utan egna anställda ingenjörer, denna byggnad  riskerar att falla samman.",
"##chatioteer_school_no_workers##":"Utan hantverkare kan inga nya vagnar produceras. Som resultat kan hippodromen, om den är i drift, bli lidande.",
"##barracks_bad_weapons_bad_workers##":"Med minimal personal och utan vapen i lager, får vi kämpa för att utbilda till och med de mest enkla trupper.",
"##fort_legionaries_no_workers##":"Utan personal kan vi inte utbilda en enda ny rekryt. Mars hjälpe oss i krigstid!",
"##militaryAcademy_no_workers##":"Utan personal kan vi inte finslipa kunskaperna för stadens nya soldater. De tvingas att gå direkt till sina poster och hoppas på det bästa.",
"##forum_no_workers##":"Utan indrivare bidrar det här kontoret inte med någonting till stadskassan.",
"##prefecture_no_workers##":"Utan personal blir den här stationen inte mycket mer än en måltavla för vandaler.",
"##tower_no_workers##":"Utan bemanning har vi ingen personal till våra katapulter eller vakter som kan patrullera murarna.",
"##gladiator_pit_no_workers##":"Utan utbildningspersonal kan denna skola inte utbilda nya gladiatorer.",
"##lion_pit_no_workers##":"Utan personal kan detta lejonhus inte leverera några nya lejon till spelen.",
"##idle_factory_in_city##":"overksam industri i staden",
"##idle_factories_in_city##":"overksamma industrier i staden",
"##wt_homeless##":"Hemlös",
"##extm_security_tlp##":"Säkerhet",
"##senatepp_unemployment##":"Arbetslöshet",
"##advchief_workless##":"Staden har en arbetslöshet på",
"##migration_lack_workless##":"Arbetslöshet minskar antalet immigranter.",
"##priest_high_workless##":"Arbetslösheten är oroväckande hög",
"##advemployer_panel_workless##":"Arbetslös arbetsstyrka ",
"##ovrn_unemployed##":"Arbetslös",
"##rioter_in_city_title##":"Vandalism i staden",
"##rioter_in_city_text##":"Vandalism i staden",
"##library##":"Bibliotek",
"##wt_librarian##":"Bibliotekarie",
"##ovrm_library##":"Bibliotek",
"##libraries##":"Bibliotek",
"##favor##":"Gynna
",
"##senatepp_favour_rating##":"Gynna
",
"##wndrt_favour##":"Gynna
",
"##thanks_to##":"TACK TILL:",
"##rome_gratitude_request_title##":"Kjesarens tacksamhet.",
"##carthago_win_text##":"Tack vare din briljanta insats ligger det karthagiska hotet äntligen bakom oss. Våra forna fiender är nu laglydiga romerska medborgare. I alla fall de som ännu är i livet!",
"##advemp_emperor_favour##":"Kjeserlig förmån
",
"##blessing_of_venus_title##":"En gudagåva från Venus",
"##spirit_of_mars_title##":"En gudagåva från Mars",
"##blessing_of_mercury_title##":"En gåva från Merkurius",
"##blessing_of_neptune_title##":"En gåva från Neptunus",
"##blessing_of_ceres_title##":"En gudagåva från Ceres",
"##romeGuard_gods_angry##":"Gudarna är rasande över denna plats!",
"##barber_gods_angry##":"Gudarna är rasande. Jag önskar att ståthållaren kunde bygga fler tempel.",
"##gods_wrathful_title##":"Gudarna är vreda",
"##doctor_gods_angry##":"Om vi inte respekterar gudarna mer, kommer vi att få känna på deras vrede.",
"##lionTamer_gods_angry##":"Gudarna är så rasande att det påverkar mitt Lejon! Han är rytande arg!",
"##legion_morale##":"Moral",
"##legion_morale_is_too_low##":"Legionens stridsmoral är för dålig för att kunna svara!",
"##rladv_mood##":"Gudarna är",
"##hospital##":"Sjukhus",
"##hospitals##":"Sjukhus",
"##big_villa##":"Stor villa",
"##big_shack##":"Stor koja",
"##big_tent##":"Stort tält",
"##statue_big##":"Stor staty",
"##big_hovel##":"Stort skjul",
"##big_hut##":"Stort hus",
"##citizens_like_chariot_races##":"Medborgarna vet inget bättre än vagnkapplöpningar.",
"##large_temples##":"Stora tempel",
"##bldm_big_temple##":"Stora tempel",
"##large##":"Stort",
"##middle_festival##":"Stor festival",
"##big_palace##":"Stort palats",
"##big_domus##":"Stor Insula",
"##large_temple##":"Stort tempel",
"##briton##":"En britt",
"##britons##":"Britter",
"##waiting_for_free_dock##":"Har kastat ankar, i väntan på ledig kajplats",
"##destroy_bridge_warning##":"Ta ned broar med försiktighet. Isolerade samhällen kommer försvinna utan tillgång till huvudvägen till Rom.
",
"##wt_rioter##":"Upprorsman",
"##no_culture_building_in_city##":"Du har ingen kultur i din stad, ergo (latin för därför!) har du ingen kulturställning.",
"##have_less_academy_in_city_0##":"Du har för få högskolor i din stad. Om du bygger fler förbättras din ställning.",
"##have_less_library_in_city_0##":"Du har för få bibliotek i din stad. Om du bygger fler förbättras din ställning.",
"##have_less_theater_in_city_0##":"Du har för få teatrar i din stad. Om du bygger fler förbättras din ställning.",
"##have_less_school_in_city_0##":"Du har för få skolor i din stad. Om du bygger fler förbättras din ställning.",
"##have_less_temple_in_city_0##":"Du har för få religiösa byggnader i din stad. Om du bygger fler förbättras din ställning.",
"##god_exalted##":"Exalterad",
"##mission_wnd_tocity##":"Till staden",
"##education_awesome##":"Alla som kräver utbildningsmöjligheter i staden har dem, och dessa är perfekta i hela staden.",
"##no_people_in_city##":"Inga människor i staden!",
"##advchief_employers_ok##":"Staden har inga arbetslöshetsproblem",
"##no_industries_in_city##":"Inga industrier i staden",
"##advchief_health_awesome##":"Stadens hälsosituation är utmärkt.",
"##advchief_health_awesome_clinic##":"Stadens hälsosituation är utmärkt, inga väntetider alls för besök till lokala läkare.",
"##city_have##":"Stadens skattkammare har tillgångar på",
"##healthadv_not_need_health_service_now##":"För närvarande finns ingen efterfrågan på hälsovård eller sanitära inrättningar. I takt med att staden utvecklas, kommer dock befolkningen att kräva badhus och sjukhus, och senare även barberare!",
"##working_have_some_labor_access##":"Denna byggnad har för närvarande viss tillgång till arbetskraft",
"##working_have_good_labor_access##":"Denna byggnad har för närvarande god tillgång till arbetskraft",
"##working_have_no_labor_access##":"Denna byggnad har för närvarande ingen tillgång till arbetskraft",
"##working_have_awesome_labor_access##":"Denna byggnad har för närvarande utmärkt tillgång till arbetskraft",
"##entadv_small_city_not_need_entert##":"För tillfället har dina medborgare andra enklare behov, än underhållning att tänka på. Men i takt med att staden växer kommer de ha begär för något som minskar enformigheten i deras vardagsliv.",
"##working_have_very_little_labor_access##":"Denna byggnad har för närvarande mycket liten tillgång till arbetskraft",
"##working_have_bad_labor_access##":"Denna byggnad har för närvarande dålig tillgång till arbetskraft",
"##its_very_peacefull_province##":"Kjesaren har aldrig förut skådat en sådan fridfull stad förut!",
"##to_empire_road##":"Till Imperiet",
"##senate_save##":"i stadskassan",
"##some_amphitheaters_no_actors##":"Vissa av dina amfiteatrar saknar skådespelare och gladiatorer. Fler underhållare skulle ge bättre villkor i de stadsdelar som klagar över dålig underhållning.",
"##advchief_high_crime_in_district##":"Vissa områden har hög kriminalitet",
"##advchief_which_crime_in_district##":"Vissa områden har mindre problem",
"##colege_access_perfectly##":"Alla områden som kräver utbildningsmöjligheter har tillgång till dem, men fler högskolor skulle minska storleken på klasserna.",
"##library_access_perfectrly##":"Alla områden som kräver utbildningsmöjligheter har tillgång till dem, men fler bibliotek skulle minska trängseln.",
"##school_access_perfectly##":"Alla områden som kräver utbildningsmöjligheter har tillgång till dem, men fler skolor skulle minska storleken på klasserna.",
"##none_crime_risk##":"Ingen brottslighet i sikte här.",
"##lost_money_last_year##":"Förra året förlorade din stad pengar - detta minskade stadens välstånd.",
"##no_food_stored_last_month##":"INGEN MAT lagrad förra månaden!",
"##to_rome_road##":"Till Rom",
"##furniture_workshop_bad_work##":"Med nästan inga snickare i verkstan, står produktionen nästan stilla. Det kommer inte att produceras mycket möbler under det kommande året.",
"##clay_pit_bad_work##":"Med nästan inga grävare vid detta lertag, står produktionen nästan helt still. Det kommer inte att produceras mycket lera under det kommande året.",
"##lumber_mill_bad_work##":"Det finns nästan inga skogsarbetare, produktionen står nästan helt still.",
"##quarry_bad_work##":"Med nästan inga anställda vid det här stenbrottet. Det kommer inte att produceras mycket marmor det kommande året.",
"##iron_mine_bad_work##":"Med nästan inga gruvarbetare här, står nästan produktionen helt still. Det kommer inte produceras mycket järn det kommande året.",
"##fruit_farm_slow_work##":"Med nästan inga anställda vid dem här fruktodlingen, kommer det ta evigheter att få någon frukt här.",
"##vegetable_farm_bad_work##":"Det finns knappt några anställda för att underhålla jordbruket, de få grönsakerna kommer att bli offer för insekter.",
"##vinard_bad_work##":"Det finns nästan inga anställda på denna vinodling. Som resultat kommer mycket få druvor att klara sig till skörden.",
"##olive_farm_bad_work##":"Med nästan inga anställda här, de flesta olivträd saknar oliver.",
"##wine_workshop_bad_work##":"Med så få anställda står produktionen nästan still. Det kommer att produceras mycket lite vin under det kommande året.",
"##oil_workshop_bad_work##":"Med nästan inga anställda i olivodlingen, har produktionen avtagit. Det kommer produceras mycket lite olivolja det kommande året.
",
"##weapons_workshop_bad_work##":"Med så få anställda står produktionen nästan still. Det kommer inte att produceras många vapen under det kommande året.",
"##pottery_workshop_bad_work##":"Med så få anställda vid krukmakeriet står produktionen nästan stilla. Det kommer inte att produceras mycket krukor under det kommande året.",
"##meat_farm_bad_work##":"Det finns knappt några anställda vid den här farmen, djurantalet e lågt och växer extremt långsamt.",
"##cartPusher_average_life##":"Flytta kärror hela dagarna är knappast kul, men att leva här gör det möjligt.",
"##sldr_terrified##":"Livrädd",
"##overall_people_are_leaving_city##":"Generellt sett, lämnar folket din stad.",
"##overall_people_are_coming_city##":"Generellt sett, kommer folket till din stad, eller vill de komma.",
"##overall_city_population_static##":"Invånarantalet i din stad är i stort sett statiskt.",
"##weapons_workshop_full_work##":"Denna smedja har alla anställda den behöver, den arbetar fullt ut med att producera vapen.",
"##furniture_workshop_full_work##":"Detta snickeri har full sysselsättning, och arbetar fullt ut med att producera möbler.",
"##pottery_workshop_full_work##":"Detta krukmakeri har alla anställda det behöver. Det arbetar fullt ut med att producera krukor.",
"##furniture_workshop_patrly_workers##":"Detta snickeri har lediga platser. Möbelproduktionen blir effektivare när de fyllts.",
"##furniture_workshop_need_some_workers##":"Detta snickeri är underbemannat, och det tar längre tid att producera möbler än vad det borde.",
"##weapons_workshop_need_some_workers##":"Denna smedja är underbemannad, och det tar längre tid att producera vapen än vad det borde.",
"##pottery_workshop_need_som_workers##":"Detta krukmakeri är underbemannat och produktionen tar längre tid än normalt.",
"##weapons_workshop_no_workers##":"Denna vapenfabrik har inga anställda. Produktionen har upphört.",
"##furniture_workshop_no_workers##":"Denna verkstad har inga anställda. Produktionen har upphört.",
"##weapons_workshop_slow_work##":"Mycket få människor arbetar i vapenfabriken. Som resultat är vapenproduktionen långsam.",
"##reservoir_info##":"Denna gigantiska cistern innehåller rent dricksvatten, som distribueras via rör av lera över en stor radie i staden. Akvedukter kan länka samman reservoarerna över stora avstånd.",
"##no_tax_in_this_year##":"Hittills i år har ingen skatt betalats från detta hus",
"##how_to_grow_prosperity##":"Ställningen har inte förändrats detta året. Att visa vinst i stadens årliga räkenskaper är det bästa sättet att förbättra välståndsställningen.",
"##citizen_low_entertainment4##":"Man kan inte roa sig alls på det här stället!",
"##prefect_so_hungry##":"Det finns inte nog med mat i staden. Det ökar brottsligheten.",
"##house_pay_tax##":"Taxbetalande hus
",
"##actor_need_workers##":"Det finns helt enkelt inte tillräckligt med arbetare i staden.",
"##house_food_only_for_month##":"Detta hus har matförråd som åtminstone kommer att räcka under den kommande månaden",
"##house_have_not_food##":"Detta hus har inget livsmedelsförråd",
"##house_have_some_food##":"Detta hus kommer snart att äta upp sitt begränsade livsmedelsförråd",
"##trouble_colloseum_no_shows##":"Detta colosseum har inga föreställningar. Det behövs gladiatorer och lejon för att locka publik.",
"##legion_haveho_soldiers_and_barracks##":"Denna legion har för närvarande inga soldater. Den existerar bara till namnet och utan förläggningar i staden kan den inte ta emot några nya trupper.",
"##legion_haveho_soldiers##":"Denna legion har för närvarande inga soldater. Den existerar bara till namnet. Endast när nyligen utbildade trupper anländer från förläggningarna kommer den att förvandlas till en stridande enhet.",
"##no_people_in_this_locality##":"Inga människor på denna plats.",
"##low_crime_risk##":"Brott inträffar sällan i detta område",
"##enemy_army_attack_city##":"En fiendes armé marserar i detta nu direkt mot dig stad. De har plundrat några städer i närheten, och de är beräknade att nå din stad detta år.",
"##weapons_workshop_need_resource##":"Denna verkstad kräver leverans av järn, från ett magasin eller från ett malmbrott, för att producera vapen.",
"##valencia_title##":"Valentia: en relativt fredlig provins",
"##low_desirability##":"Du behöver göra området mer attraktivt -kanske genom att anlägga några trädgårdar eller torg.",
"##wn_barbarian##":"Barbar",
"##barbarian_attack_title##":"Barbarer anfaller!",
"##cant_calc_prosperity##":"Din stad är ny. Vi har inte haft möjlighet att bedöma ditt välstånd än!",
"##big_fest_description##":"Din 2 dagars festival för din valda gud är slut. Ditt folk respekterar dig.",
"##governor_palace_1_info##":"Ditt hem är en av stadens mest attraktiva adresser.",
"##not_enought_place_for_legion##":"Din legion har de fort som krävs",
"##playerarmy_gone_to_home##":"Din legion på återtåg till din stad",
"##playerarmy_gone_to_location##":"Din legion marscherar för att befria en stad från riket",
"##trade_advisor_blocked_wine_production##":"Din handelsrådgivare har stoppat all vinproduktion.",
"##trade_advisor_blocked_oil_production##":"Din handelsrådgivare har stoppat all oljeproduktion.",
"##trade_advisor_blocked_furniture_production##":"Din handelsrådgivare har stoppat all möbeltillverkning.",
"##trade_advisor_blocked_weapon_production##":"Din handelsrådgivare har stoppat all vapenproduktion.",
"##trade_advisor_blocked_grape_production##":"Din handelsrådgivare har stoppat all druvodling.",
"##trade_advisor_blocked_vegetable_production##":"Din handelsrådgivare har stoppat all grönsaksodling.",
"##trade_advisor_blocked_olive_production##":"Din handelsrådgivare har stoppat all olivodling.",
"##trade_advisor_blocked_wheat_production##":"Din handelsrådgivare har stoppat all veteodling.",
"##trade_advisor_blocked_meat_production##":"Din handelsrådgivare har stoppat all köttproduktion.",
"##trade_advisor_blocked_fruit_production##":"Din handelsrådgivare har stoppat all fruktodling.",
"##trade_advisor_blocked_timber_production##":"Din handelsrådgivare har stoppat all avverkning.",
"##trade_advisor_blocked_clay_production##":"Din handelsrådgivare har stoppat alla lertag.",
"##trade_advisor_blocked_marble_production##":"Din handelsrådgivare har stoppat all marmorbrytning.",
"##trade_advisor_blocked_iron_production##":"Din handelsrådgivare har stoppat all malmbrytning.",
"##trade_advisor_blocked_pottery_production##":"Din handelsrådgivare har stoppat all kruktillverkning.",
"##your_salary_frowned_senate##":"I Rom ser man ner på din fräckhet att betala dig själv en lön som är högre än din rang.",
"##broke_empiretax_warning##":"Din oförmåga att betala tribut till Rom utmålar din stad som misslyckad.",
"##broke_empiretax_with2years_warning##":"Din fortsatta oförmåga att lämna tribut till Rom skadar ditt rykte.",
"##your_favour_increased_from_last_year##":"Din ställning i Rom har förbättrats sedan förra året.",
"##your_favour_unchanged_from_last_year##":"Din ställning är oförändrad sedan förra året.",
"##lugdunum_win_text##":"Din behandling av gallerna i Lugdunum och den sköna stadens prakt bådar väl för Roms expansion i den norra vildmarken. Bra gjort!",
"##capua_win_text##":"Din förmåga att styra imponerar på mig. Många ståthållares karriärer gäckas när jag ber dem bygga den första kolonin. Ledare som du garanterar Rom en framtid. Kan du upprepa dina framgångar eller var det bara tur?",
"##city_need_workers_text##":"Din stad behöver fler arbetare
",
"##city_need_more_workers##":"Din stad kräver fler arbetare",
"##more_0_month_from_festival##":"Ditt folk, somliga fortfarande berusade efter festen, välkomnar din generositet.",
"##desirability_indiffirent_area##":"Dina medborgare ser varken positivt eller negativt på detta område",
"##more_12_month_from_festival##":"Ditt invånare är mycket missnöjda med tanken på ännu ett år utan en festival.",
"##need_temples_for_city##":"Dina medborgare har börjat bli intresserade av religion. Frånvaron av en närliggande gudstjänstplats hindrar stadens utveckling.",
"##gods_unhappy_text##":"Dina medborgarna tror att gudarna kan bli upprörda. Vissa medborgare har visioner av annalkande katastrofer. Bygg nya tempel och börja fester för deras skull, annars riskerar du att drabbas av deras vrede.",
"##small_colloseum_show##":"Det krävs fler spektakel i dina colosseum! Genom att förse dem med gladiatorer eller lejon förbättras underhållningen i delar av staden.",
"##send_legion_to_emperor##":"Be din militära rådgivare att avdela några stridsklara legioner i imperiets tjänst",
"##venus##":"Venus",
"##smcurse2_of_venus_description##":"Venus kastar en svart skugga av förtvivlan över din stad, vilket sätter ner humöret på dina vanvördiga medborgare.",
"##smcurse_of_venus_title##":"Venus är upprörd",
"##blessing_of_venus_description##":"Venus förmedlar en känsla av välvilja till din stad, vilket får alla dina medborgare på bättre humör.",
"##smcurse_of_venus_description##":"Venus, förmedlare av kärlek och harmoni, är upprörd. Detta bådar inget gott för prefekterna i din stad!",
"##return_2_fort##":"Återvänd till fortet",
"##return_to_main_map##":"Återvänd till spelets huvudkarta",
"##shipyard##":"Fartygsvarv",
"##wt_romeHorseman##":"Beridna stödtrupper",
"##wn_visigoth##":"Visigoter",
"##city_loathed_you##":"Du föraktas i hela staden",
"##explosion##":"Explosion",
"##varieties_food_eaten##":"Olika sorters livsmedel som ätits,",
"##governor_palace_2##":"Ståthållarens villa",
"##governorVilla##":"Ståthållarens villa",
"##wine##":"Vin",
"##prettyWine##":"Falern Vin",
"##grape##":"Vindruvor",
"##vinard_info##":"Druvorna från dessa vinrankor har odlats särskild för vinframställning. Vingårdarna gör fint vin för dina egna patricier, samt för export.",
"##vinard##":"Druvodling",
"##wine_workshop_info##":"Vinhandlare förvandlar druvor till vin, vilket patricierna kräver om de skall bygga villor. Vin är en handelsvara som är begärlig för många.",
"##wine_workshop##":"Vingård",
"##tradeadv_industrystate_tip##":"Starta eller avsluta produktion för denna aktivitet överallt i staden",
"##city_opts_god_on##":"Gudar: På",
"##city_opts_god_off##":"Gudar: Av",
"##warning##":"Varningar",
"##warehouse_gettinfull_warning##":"VARNING Denna lagerbyggnad håller på att bli full. Den kan bara ta emot varor som redan finns, inga nya varutyper.",
"##warehouse_full_warning##":"VARNING Denna lagerbyggnad är helt fylld. Den kan inte ta emot fler varor.",
"##changesalary_greater_salary##":"Varning: Betala dig själv en lön som överstiger din grad imponerar inte på kejsaren.",
"##working_build_poor_labor_warning##":"Varning: Dålig tillgång till arbetskraft",
"##working_building_need_road##":"VARNING. Denna byggnad fungerar ej. Den ligger inte intill en väg, och dess anställda kommer ej fram",
"##ovrm_water##":"Vatten",
"##water_caption##":"Vatten",
"##massilia_preview_mission##":"Det enda vattnet finns i oasen. Detsamma gäller tyvärr för odlingsbar mark. Reservoarer och lantgårdar konkurrerar om samma utrymme. Använd det med förstånd.",
"##water_info##":"Kan inte forceras, men broar kan byggas på vissa platser. Vatten är en vital handelslänk till resten av imperiet via handelshamnar. Lertag måste byggas nära vatten.",
"##water_supply##":"Vatten",
"##militaryAcademy##":"Militärhögskola",
"##advchief_military##":"Militär",
"##adve_military##":"Militär",
"##high_salary_angers_senate##":"Den löjligt höga lön du betalar till dig själv upprör senaten. Hela Rom talar om din öppna girighet.",
"##charioteer##":"Körsven",
"##citychart_census##":"Folkräkning",
"##wn_helveti_soldier##":"En helvetisk soldat",
"##barbarian_warrior##":"En barbarisk soldat",
"##wn_visigoth_soldier##":"En visigotisk soldat",
"##wn_gaul_soldier##":"En gallisk soldat",
"##goth_warrior##":"En gotisk soldat",
"##hun_warrior##":"En hunnersoldat",
"##wn_celt_soldier##":"En keltisk soldat",
"##wt_pict_soldier##":"En piktisk soldat",
"##mars_desc##":"Krig",
"##migration_war_deterring##":"Krig avskräcker immigranter!!",
"##RomeChastenerArmy_troops_at_our_gates##":"Imperiets trupper står vid stadsportarna",
"##wt_wolf##":"Varg",
"##lgn_wolves##":"Vargarna",
"##request_failed##":"Din nyligen visade oförmåga eller ovilja att utföra en kejserlig begäran har skadat din ställning i Rom en aning.",
"##market_kid_say_1##":"Den tjocka damen bad mig bära detta och följa efter henne.",
"##sldr_encouraged##":"Uppmuntrad",
"##gatehouse##":"Grindstuga",
"##more_8_month_from_festival##
":"Minnet av den tidigare festivalen håller på att blekna.",
"##east##":"Öst",
"##delighted##":"Förtjusta",
"##lionTamer_average_life##":"Här är lite utländskt kött åt dig, Leo.",
"##100_citizens_in_city##":"Din stads population har nått 100 invånare för första gången.",
"##1000_citizens_in_city##":"Din stads population har nått 1.000 invånare för första gången.",
"##10000_citizens_in_city##":"Din stads population har nått 10.000 invånare för första gången.",
"##15000_citizens_in_city##":"Din stads population har nått 15.000 invånare för första gången.",
"##2000_citizens_in_city##":"Din stads population har nått 2.000 invånare för första gången.",
"##20000_citizens_in_city##":"Din stads population har nått 20.000 invånare för första gången.",
"##25000_citizens_in_city##":"Din stads population har nått 25.000 invånare för första gången.",
"##3000_citizens_in_city##":"Din stads population har nått 3.000 invånare för första gången.",
"##500_citizens_in_city##":"Din stads population har nått 500 invånare för första gången.",
"##5000_citizens_inc_city##":"Din stads population har nått 5.000 invånare för första gången.",
"##enemies_attack_title##":"Fiender attackerar staden",
"##city_have_defence##":"Stadens försvar skulle aldrig ha släppt igenom fienden!",
"##enemies_at_the_door##":"Fiender vid dina portar",
"##barbarian_are_closing_city##":"Fiender närmar sig staden",
"##barbarian_attack_text##":"Roms fiender är i utkanten av din stad. Räkna med 1 flaska vin eller 2 - och vad de mer önskar sig.",
"##enemy_army_threating_a_city##":"En fiendearmé som hotar en av rikets städer",
"##city_under_barbarian_attack##":"Fiendesoldaterna i stadens omgivning förbättrar inte din fredsställning!",
"##time_since_last_gift##":"Tid sedan senaste gåva",
"##ovrm_education##":"Allt",
"##ovrm_entertainment##":"Allt",
"##religionadv_need_basic_religion##":"Fler och fler medborgare kräver minst en gudstjänstplats i sitt bostadsområde, för att förbättra gudarnas uppfattning om dem.",
"##healthadv_some_regions_need_doctors_2##":"Fler och fler människor vill ha bekväm tillgång till hälsovård. Anordna lokal tillgång till kliniker så att staden kan växa.",
"##for_second_year_broke_tribute##":"För andra året i rad har du inte betalat tribut till Rom. Detta håller på att bli ett stort problem för din framtida karriär.",
"##tarsus_win_text##":"Du är på god väg att bli min mest uppskattade undersåte. Din mästerliga förståelse av handeln gjorde Tarsus till precis den stad jag hoppats på. De östliga provinserna är mer lojala i dag, tack vare dig.",
"##tutorial2_win_text##":"Du lär dig snabbt! Nu har du tillräckligt med kunskap för att klara ett riktigt uppdrag. Från och med nu kan du välja vilken riktning din karriär ska ta. Välj en fredligare provins om du vill koncentrera dig på att styra eller en farligare provins om du vill tampas med Roms fiender.",
"##taxCollector_high_tax##":"Har du sett skatterna här? Medborgare, det är inte rätt.",
"##can_build_only_one_of_building##":"Du kan endast ha en byggnad av denna typ",
"##emperor_anger_text##":"Du avsikligt vägrar skicka mig det jag frågat efter? Eller vill du förnedra mig?",
"##imperial_reminder_text##":"Har du glömt bort min senaste förfrågan? Jag börjar tappa tålamodet.",
"##emigrant_high_workless##":"Vet ni var det kan finnas arbete? Jag måste få ett arbete.",
"##current_year_notpay_tribute_warning##":"Du har inte betalat tribut detta året. Spara lite pengar i din skattkammare så att du kan göra din årliga betalning.",
"##request_faild_text#":"Du trotsar mig fortfarande? Strunta i min förfrågan. Jag söker någon annanstans. Du ska ha tur om jag återvänder.",
"##ive_asked_senate_proclaim_you_a_god##":"Gratulerar! Du har uppnått de högsta poängställningar som någonsin åstadkommits av Roms ståthållare. Jag är stolt över att få lämna över till dig. Jag kungör att du må krönas till kejsare och härskare över hela imperiet. Äntligen kan jag dra mig tillbaka till min villa på ön, som en vanlig medborgare igen. Må ditt namn...",
"##wrath_of_neptune_failed_description##":"Du har åtdragit mitt vrede. Jag ser fram emot när din stad börjar använda båtar, då kommer hämnden.",
"##sentiment_people_annoyed_you##":"Människorna är irriterade på dig",
"##city_has_runout_money_again##":"Du har slösat med Roms tillgångar. Caesar har ilsket gått med på att låna 5.000 denarii for 12 månader. Du behöver generera pengar från skatt och exportering.",
"##damascus_win_text##":"Ännu en gång har du uppnått vad svagare män kallar omöjligt. Hela östern åsåg din balansgång i Damaskus. Nu kan jag tryggt hämta hem några av mina syriska legioner.",
"##really_destroy_fort##":"Är du säker på att du vill ta detta fort ur aktiv tjänst?",
"##tingis_win_text##":"Är du ståthållare eller general? Din utmärkta insats vid Tingis befriar mina legioner från tjänstgöring i väst och låter mig ägna tiden åt andra strävanden. Du börjar bli en nyckelperson i min planering.",
"##enter_your_name##":"Välj ett namn",
"##select_location##":"Välj destination",
"##select_city_layer##":"Välj en översiktsrapport för staden",
"##priority_button_tolltip##":"Klicka på ett nummer för att fastställa prioritetsnivå. Alla övriga uppgifter kommer att omjusteras",
"##select_this_graph##":"Välj detta diagram",
"##mainmenu_language##":"Språk",
"##exit_without_saving_question##":"Avsluta utan att spara?",
"##gmenu_file_mainmenu##":"Avsluta till huvudmenyn",
"##gmenu_exit_game##":"Avsluta spel",
"##gmenu_file_exit##":"Avsluta spel",
"##mainmenu_quit##":"Avsluta spel",
"##exit_salary_window##":"Lämna löneskärmen",
"##donationwnd_exit_tip##":"Lämna donationsskärmen",
"##exit_this_panel##":"Avsluta denna panel",
"##migration_broke_workless##":"Hög arbetslöshet i din stad bromsar din välståndsställning.",
"##migration_broke_tax##":"Höga skatter gör att vissa människor undviker din stad",
"##migration_middle_lack_tax##":"Höga skatter förhindrar immigration",
"##high_fire_risk##":"Stor brandrisk",
"##high_damage_risk##":"Stor risk att kollapsa",
"##migration_lack_crime##":"Hög brottslighet skrämmer lokalbefolkningen.",
"##quit##":"Avsluta",
"##exit##":"Avsluta",
"##wn_gaul##":"Galler",
"##egift_gaulish_bodyguards##":"Galliska livvakter",
"##egift_gepards_and_giraffes##":"Geparder och giraffer",
"##lgn_heroes##":"Hjältarna",
"##lgn_hydras##":"Hydrorna",
"##chief_advisor##":"Huvudrådgivare",
"##wt_gladiator##":"Gladiator",
"##gladiator_bouts_runs_for_another##":"Gladiatorkampen pågår ytterligare",
"##amphitheater_haveno_gladiator_bouts##":"Ingen gladiatorkamp för närvarande",
"##colloseum_haveno_gladiator_bouts##":"Ingen aktuell gladiatorkamp",
"##clay##":"Lera",
"##clay_pit##":"Lertag",
"##gods_unhappy_title##":"Gudar är missnöjda",
"##wrath_of_venus_title##":"Venus vrede",
"##emperor_anger##":"Kjesarens ilska",
"##wrath_of_mars_title##":"Mars vrede",
"##smallcurse_of_mars_failed_title##":"Mars vrede",
"##wrath_of_mercury_title##":"Mercury vrede",
"##wrath_of_neptune_title##":"Neptune vrede",
"##wrath_of_ceres_title##":"Ceres vrede",
"##immigrant_much_food_here##":"De påstår att det finns mat här. Är det en bra plats att bo på?",
"##year##":"Sädesmagasin lagrar",
"##charioter_so_hungry##":"Hungrig? Jag kan äta en häst, så lite mat finns det.",
"##hippodrome_haveno_races##":"Inga kapplöpningar för närvarande",
"##current_races_runs_for_another##":"Kapplöpningar pågår ytterligare",
"##pottery_workshop##":"Krukmakeri",
"##city##":"Stad",
"##city_in_debt##":"Stad i skuld",
"##city_fire_title##":"Eldsvåda i din stad",
"##city_still_in_debt##":"Stad fortfarande i skuld",
"##pestilent_event_text##":"En farsot har drabbat staden. Bristen på sjukhus fordrar att dina prefekter desinfekterar de drabbade stadsdelarna.",
"##city_is_besieged##":"Staden är belägrad",
"##city_in_debt_again##":"Stad i skuld igen",
"##city_health##":"Hälsosituation",
"##city_sounds_on##":"Stadsljud är på",
"##city_sounds_off##":"Stadsljud är av",
"##advchief_needworkers##":"Staden saknar",
"##citizens_enjoy_drama_and_comedy##":"Medborgarna njuter av drama och komedi enligt den grekiska traditionen.",
"##citizens_here_are_bored_for_chariot_races##":"Medborgarna är uttråkade. Trots hästkapplöpningarna finns det inte tillräckligt med underhållning här.",
"##burning_ruins##":"Brinnande ruin",
"##ovrm_hospital##":"Sjukhus",
"##wn_goth##":"Gother",
"##not_need_education##":"Inga medborgare kräver ännu utbildningsmöjligheter. Men när staden börjar växa kommer människor att förvänta sig skolor och högskolor, och senare även bibliotek.",
"##gods_wrathful_text##":"Medborgarna fruktar att minst en av gudarna hyser vrede mot staden. De bönfaller dig att bygga fler tempel för att blidka dem.",
"##citizen_are_rioting##":"Medborgarna gör uppror!",
"##doctor_good_life##":"Stadens invånare tycks vara vid god hälsa.",
"##well_info##":"Medborgare utan tillgång till fontän kan ta vatten från brunnar, men stadsdelar med brunnsvatten är inga trevliga platser att bo på.",
"##patrician_gods_angry##":"Medborgare! Situationen är hotfull. Gudarna är vreda.",
"##patrician_low_entertainment##":"Medborgare! Är icke detta den tråkigaste staden i riket?",
"##recruter_need_workers##":"Medborgare! Denna stad behöver fler arbetare.",
"##gladiator_perfect_life##":"Medborgare! Jag har kämpat i många städer och den här är en av de bästa.",
"##citizen##":"Medborgare",
"##great_festival##":"Storslagen festival",
"##mopup_formation_title##":"Upprensningsformation",
"##wn_graeci##":"Greker",
"##egift_gree_manuscript##":"Ett grekiskt manuskript",
"##greek_soldier##":"En grekisk soldat",
"##gmsndwnd_game_volume##":"Volym",
"##yes##":"Ja",
"##citizen_low_salary##":"Min hund skulle inte arbeta för de löner de betalar här. Jag ger mig av.",
"##city_damascus##":"Damascus",
"##damascus_title##":"Damaskus: en relativt farlig provins",
"##donation_is##":"Donationen är",
"##date_tooltip##":"Datum",
"##date##":"Datum",
"##scrw_date##":"Datum",
"##governor_palace_3##":"Ståthållarens palats",
"##governorPalace##":"Ståthållarens palats",
"##month_12_short##":"Dec",
"##dn's##":"Avsluta byggare",
"##dn_per_month##":"denarer per månad",
"##dn_collected_this_year##":"denarer har betalats hittills i år",
"##dn##":"Spara karta",
"##day##":"Dag",
"##funds_tooltip##":"Kassa",
"##trees_and_forest_caption##":"Träd och skogsland",
"##children##":"Barn",
"##srcw_no_messages##":"Inga nya meddelanden",
"##need_barracks_for_work##":"Fungerande förläggning krävs för att ta emot soldater",
"##tower_need_wall_for_patrol##":"Måste finnas intill en mur för att sända ut en patrull",
"##need_marble_for_large_temple##":"Du behöver 2 ton marmor för att bygga ett stort tempel",
"##oracle_need_2_cart_marble##":"Du behöver 2 ton marmor för att bygga ett orakel",
"##furniture_workshop_need_resource##":"Detta snickeri behöver leverans av virke från ett magasin eller från en brädgård för att kunna producera möbler.",
"##pottery_workshop_need_resource##":"Detta krukmakeri behöver leveranser av lera, från ett magasin eller från ett lertag, för att kunna producera krukor.",
"##need_access_to_full_reservoir##":"Kräver tillgång till en full reservoar för att fungera",
"##haveno_trade_routes_for_goods##":"Det finns inga öppna handelsvägar för dessa varor",
"##advemployer_panel_denaries##":"dn",
"##denarii_short##":"dn",
"##days##":"Dagar",
"##age_bc##":"BC",
"##bc##":"fKr",
"##marketBuyer_good_life##":"God dag, medborgare. Är det inte en härlig stad?",
"##clay_pit_info##":"Tag lera och handla med, eller leverera den till krukmakerier. Folket behöver krukor för att bebo Insulaen.",
"##iron_mine_info##":"Bryt järn för att handla med, eller för att leverera till vapensmedjorna. Utrusta din armé med hemgjorda vapen, eller exportera dem till andra provinser.",
"##quarry_info##":"Bryt marmor ur intilliggande klippor och använd den till att bygga orakel och stora tempel. Marmor är vanligen en värdefull exportvara.",
"##god_pleased##":"Nöjda",
"##sld_quite_daring##":"Mycket djärv",
"##blessing_of_neptune_description##":"Glad över ditt växande intresse för honom garanterar Neptunus alla dina sjöfarande handelsmän lugna seglatser under resten av året. De kommer att betala dig dubbelt under den tiden.",
"##dock##":"Handelshamn",
"##wt_docker##":"Hamnarbetare",
"##ovrm_clinic##":"Kliniker",
"##clinic_info##":"Läkares förbättrar medborgarnas hälsa genom sina hembesök i de stadsdelar som ingår i deras runda. Blomstrande områden vill ha en klinik.",
"##city_has_debt##":"Staden har en skuld till Rom på",
"##lutetia_win_text##":"Kejsar Augustus måste ha anat ditt styre när han förutspådde vår seger över gallerna. Din framgång vid Lutetia räcker långt när det gäller att krossa deras upprorsanda.",
"##marketBuyer_low_entertainment##":"Detta måste vara den tråkigaste staden i imperiet.",
"##governor_palace_1##":"Ståthållarens hus",
"##governorHouse##":"Ståthållarens hus",
"##houseBtnTooltip##":"Hus",
"##mainmenu_package##":"Advancerade inställningar",
"##package_options##":"Avancerade inställningar",
"##graphics##":"GRAFIK:",
"##advanced_houseinfo##":"Avancerad information om detta hus",
"##citizens_additional_rooms_for##":"Extra utrymme för",
"##road_caption##":"Väg",
"##road_text##":"Vägarna är livsviktiga för stadens funktion. Invånarna går bara ut ur sina hus om det finns en väg.",
"##citychart_society##":"Samhälle",
"##bath_access##":"Badtillgång",
"##barber_access##":"Barberartillgång",
"##ovrm_market##":"Marknadstillgång",
"##formation_available_for_trained_troops##
":"Endast tillgänglig för trupper som utbildats på militärhögskola.",
"##debet##":"Inkomst",
"##timber##":"Timmer",
"##spirit_of_mars_text##":"Andan väktare trollade av Mars för att skydda dig vaknar, och lägger låg några av dem som vågar angripa hans valda staden.",
"##wn_eygptian_soldier##":"En egyptisk soldat",
"##egift_egyptian_glassware##":"Egyptiska glasvaror",
"##wn_eygptians##":"Eygptier",
"##ovrm_food##":"Mat",
"##units##":"Enheter",
"##unit##":"Enhet",
"##gmspdwnd_autosave_interval##":"Spara automatiskt",
"##warning_theater_access##":"Detta hus har inte passerats av en skådespelare på ett tag. Det kommer snart att förlora tillgången till teater",
"##warning_baths_access##":"Om ingen badhusarbetare passerar snart, kommer detta hus att förlora sin tillgång till badhus",
"##warning_library_access##":"Om ingen bibliotekarie passerar huset snart, kommer det att förlora sin tillgång till bibliotek",
"##taxCollector_low_entertainment##":"Jag skulle inte ha nåt emot att pressa folk på denarer hela dagarna om det bara fanns mer att göra på kvällarna!",
"##romeGuard_low_entertainment##":"Om det fanns bättre underhållning i staden skulle vakttjänsten inte kännas så betungande.",
"##seamerchant_noany_trade##":"Om jag fick bestämma skulle jag inte segla den här vägen. Den här staden varken köper eller säljer något.",
"##lionTamer_so_hungry##":"Om vi inte får mer mat snart, äter lejonet upp mig!",
"##engineer_so_hungry##":"Om jag inte får mat snart ger jag mig av från staden.",
"##taxCollector_so_hungry##":"Om vi inte får mer livsmedel finns det snart ingen som kan betala skatt!",
"##warning_doctor_access##":"Om ingen läkare passerar huset snart, kommer det att förlora sin tillgång till läkarklinik",
"##tamer_normal_life##":"Om du rör mitt lejon, får du smaka på min piska.",
"##taxCollector_gods_angry##":"Om vi inte bygger fler tempel snart, kommer gudarna att förbanna denna stad.",
"##teacher_gods_angry##":"Vi får känna gudarnas vrede om vi inte bygger fler tempel snart.",
"##warning_barber_access##":"Om ingen barberare går förbi huset snart, kommer det att förlora sin tillgång till barberare",
"##this_fire_can_spread##":"Dessa eldsvådor sprider sig om du inte snabbt hejdar dem.",
"##warning_college_access##":"Om ingen lärare passerar huset snart, kommer det att förlora sin tillgång till högskola",
"##warning_hospital_access##":"Om ingen kirurg passerar detta hus snart, kommer det att förlora sin tillgång till sjukhus",
"##rioter_say_3##":"Om du vill veta hur städer ser ut när de brinner, se noga på nu!",
"##warning_school_access##":"Om inget skolbarn passerar huset snart, kommer det att förlora sin tillgång till skola",
"##citizen_high_workless2##":"Om jag inte får arbete snart, måste jag flytta till en annan stad.",
"##immigrant_so_hungry##":"Om jag stannar längre dör jag. Det finns ingen mat någonstans.",
"##day_longer_in_that_tent##":"En dag till i det tältet och jag hade exploderat",
"##seamrchant_another_successful_voyage##":"Ännu en lyckosam resa. Förtjänsten från denna stad gör att man står ut med sjösjukan.",
"##architect_salary##":"Arkitektlön på",
"##citizen_salary##":"Medborgarlön på",
"##engineer_salary##":"Ingenjörslön på",
"##quaestor_salary##":"Kvestorslön på",
"##clerk_salary##":"Bokhållarlön på",
"##consul_salary##":"Konsulslön på",
"##praetor_salary##":"Pretorslön på",
"##proconsoul_salary##":"Prokonsulslön på",
"##procurator_salary##":"Prokuratorslön på",
"##caesar_salary##":"Caesars lön på",
"##edil_salary##":"Edillön på",
"##more_salary_dispeasure_senate##":"Den lön som du betalar dig själv, och som vida överskrider din rang, är en källa till missnöje i Rom.",
"##prefect_fight_fire##":"Hettan från elden är otroligt stark.",
"##iron_mine##":"Malmbrott",
"##iron##":"Järn",
"##lgn_stallion##":"Hingstarna",
"##meat_farm##":"Svinuppfödning",
"##priest_good_life##":"Livet är mycket behagligt i denna stad.",
"##actor_average_life##":"Livet här är helt enkelt ljuvligt.",
"##barber_average_life##":"Är inte den här staden ett riktigt klipp?",
"##occupants##":"invånare",
"##money_stolen_title##":"Folket är arga",
"##sentiment_people_pleased_you##":"Människorna är nöjda med dig",
"##sentiment_people_extr_pleased_you##":"Människorna är extremt nöjda med dig",
"##house_not_report_about_crimes##":"De boende har inte rapporterat någon brottslighet.",
"##sentiment_people_upset_you##":"Människorna är upprörda över dig",
"##sentiment_people_love_you##":"Människorna älskar dig",
"##sentiment_people_verypleased_you##":"Människorna är mycket nöjda med dig",
"##sentiment_people_veryupset_you##":"Människorna är mycket upprörda över dig",
"##sentiment_people_veryangry_you##":"Människorna är mycket arga på dig",
"##house_provide_food_themselves##":"Tältboende hämtar sin egen mat från omgivande marker.",
"##fountain_info##":"Människorna hämtar allt vatten som de behöver från fontäner, som måste förses med vatten via ledningar från en reservoar. Fontäner är den källa till vatten som folket föredrar.",
"##sentiment_people_idolize_you##":"Människorna avgudar dig, som en gud",
"##sentiment_people_indiffirent_you##":"Människorna är likgiltiga inför dig",
"##sentiment_people_angry_you##":"Människorna är arga på dig",
"##wt_priest##":"Präst",
"##hlth_care_of##":"Sköter om",
"##load_this_game##":"Ladda",
"##mainmenu_load##":"Ladda spel",
"##mainmenu_loadgame##":"Ladda spel",
"##mainmenu_loadcampaign##":"Ladda kampanj",
"##mainmenu_loadmap##":"Ny karta",
"##Load_save##":"Öppna sparat spel",
"##mainmenu_playmission##":"Ladda scenario",
"##fileload_load_tlp##":"Öppna detta sparade spel",
"##initialize_animations##":"Laddar animationer",
"##initialize_names##":"Laddar medborgarnamnen",
"##initialize_walkers##":"Laddar fotgängarinställningar",
"##initialize_constructions##":"Laddar konstruktionsinställningar",
"##initialize_religion##":"Laddar religioninställningar",
"##loading_offsets##":"Laddar texturer",
"##initialize_house_specification##":"Laddar husdata",
"##meat_farm_info##":"Välmående medborgare njuter av olika sorters fläsk. Kött kan förvaras i sädesmagasin för lokal konsumtion eller i handelsmagasin för export.",
"##close##":"Stäng",
"##infobox_tooltip_exit##":"Stäng detta fönster",
"##wt_marketBuyer##":"Marknadsbesökare",
"##advchief_employment##":"Arbete",
"##west##":"Väst",
"##grape_factory_stock##":"Lagrade druvor,",
"##clay_factory_stock##":"Lagrad lera,",
"##timber_factory_stock##":"Lagrat virke,",
"##iron_factory_stock##":"Lagrat järn,",
"##olive_factory_stock##":"Lagrade oliver,",
"##weapon_store_of##":"Vapenupplaget har",
"##advchief_food_stocks##":"Matförråd",
"##have_food_for##":"Livsmedelsförråd för",
"##mainmenu_dlc_articles##":"Artiklar",
"##pay_to_open_trade_route?##":"Betala för att öppna denna väg?",
"##emp_pay_open_this_route_question##":"Betala för att öppna denna väg?",
"##contaminted_water##":"Förorenat vatten",
"##advemployer_panel_salary##":"Löner",
"##wages##":"Löner",
"##captured_city##":"En erövrad stad",
"##collapsed_building_title##":"Kollapsad byggnad",
"##destroyed_building_title##":"Förstörd byggnad",
"##pottery_workshop_info##":"Här formar krukmakare lera till kärl som medborgarna använder till förvaring. Handla med krukor, eller låt dina marknader distribuera dem så att människorna kan bygga bättre hus.",
"##barber_need_workers##":"Det saknas många arbetare här.",
"##some_crime_risk##":"Området löper viss risk att drabbas av brottslighet.",
"##nativeHut_info##":"En del lokalbefolkning bor här, de lever ett stillsamt enkelt liv. De vill bara bli lämnade ifred.",
"##lionTamer_high_workless##":"Det är stor arbetslöshet här.",
"##marketBuyer_so_hungry##":"Det finns inte tillräckligt med livsmedel här. Hur ska jag kunna försörja mig?",
"##teacher_so_hungry##":"Det saknas livsmedel här. Det gör medborgarna olyckliga.",
"##high_crime_risk##":"Detta område står i begrepp att explodera i upplopp.",
"##landmerchart_noany_trade2##":"Inget att byteshandla med här, passerar bara",
"##oil_workshop_info##":"Här pressas olja från oliver, som plebejerna behöver för matlagning och för belysningen i sin Insulae. Överskottsoljan kan bli lönsam handel.",
"##wheat_farm_bad_work##":"Det finns mycket få jordbruksarbetare här. Som resultat är veteproduktionen långsam.",
"##furniture_workshop_slow_work##":"Mycket få snickare arbetar här. Som resultat är möbelproduktionen långsam.",
"##olive_farm_slow_work##":"Det finns mycket få människor som arbetar här. Som resultat är olivproduktionen långsam.",
"##pottery_bad_work##":"Mycket få människor arbetar här. Som resultat går krukproduktionen långsamt.",
"##vegetable_farm_slow_work##":"Mycket få jordbrukare arbetar här. De få grönsaker som odlas är små och osunda.",
"##fig_farm_bad_work##":"Mycket få människor arbetar i denna fruktträdgård. Fruktskörden kommer att bli liten och sen.",
"##advchief_low_crime##":"Det finns lite brottslighet här, ingenting allvarligt.",
"##scholar_need_workers##":"Det finns så få arbetare att någon till och med erbjöd mig jobb.",
"##gladiator_high_workless##":"De arbetslösa är så många här. Jag önskar vi kunde få träna oss på några av dem.",
"##scholar_high_workless##":"Det är jättemånga som söker arbete här.",
"##barber_high_workless##":"Arbetslösheten är så hög att den får håret att stå på ända!",
"##actor_high_workless##":"Det är så stor arbetslöshet att jag inte förmår lära mig mina repliker.",
"##library_info##":"Litterära arbeten från hela riket förvaras här på grekiska och latin. Lärda män insisterar att biblioteken är avgörande för en viktig stad.",
"##romeGuard_average_life##":"Allt verkar lugnt här.",
"##advchief_health##":"Hälsa",
"##health##":"Hälsa",
"##ovrm_healthAll##":"Hälsa",
"##ovrm_health##":"Hälsa",
"##advchief_health_low##":"Stadens hälsosituation är förfärande",
"##advchief_health_lower##":"Stadens hälsosituation är förfärande, pest kommer med all säkerhet bryta ut.",
"##advchief_health_high##":"Stadens hälsosituation är bra",
"##advchief_health_high_clinic##":"Stadens hälsosituation är bra, dina medborgare lider bara av enklare sjukdomar.",
"##advchief_health_middle##":"Stadens hälsosituation är tillfredsställande",
"##advchief_health_middle_clinic##":"Stadens hälsosituation är tillfredsställande, klinikerna håller farliga epidemier borta.",
"##advchief_health_verygood##":"Stadens hälsosituation är mycket bra",
"##advchief_health_verygood_clinic##":"Stadens hälsosituation är mycket bra, medborgarnas småkrämpor hanteras snabbt av lokala läkare.",
"##advchief_health_less##":"Stadens hälsosituation är ganska dålig",
"##advchief_health_less_clinic##":"Stadens hälsosituation är dålig, mat och kliniker skulle förbättra hälsan.",
"##advchief_health_good##":"Stadens hälsosituation är nästan perfekt",
"##advchief_health_good_clinic##":"Stadens hälsosituation är nästan perfekt, läkarnas kliniker är nästan tomma.",
"##advchief_health_perfect##":"Stadens hälsosituation är perfekt",
"##advchief_health_perfect_clinic##":"Stadens hälsosituation är perfekt, dina tomma kliniker utgör ett exempel genom hela imperiet.",
"##advchief_health_terrible_clinic##":"Stadens hälsosituation är fruktansvärd, klinikerna hinner inte med, sjukdomar är nästan oundvikliga.",
"##advchief_health_terrible##":"Stadens hälsosituation är fruktansvärd",
"##adve_health_education##":"Hälsa och utbildning",
"##soldiers_health##":"Soldaternas hälsa",
"##extm_health_tlp##":"Hälsa",
"##ceres_desc##":"Jordbruk",
"##earthquake_title##":"Jordbävning",
"##wheat##":"Vete",
"##wheat_farm_info##":"Vetekorn är det grundläggande livsmedlet för ditt folk. Det måste lagras i sädesmagasin för att livnära ditt folk, eller i handelsmagasin för export.",
"##angry##":"Arga",
"##lgn_snakes##":"Ormarna",
"##egift_golden_chariot##":"En gyllene vagn",
"##wn_iberian_soldier##":"En iberisk soldat",
"##developers##":"UTVECKLARE:",
"##testers##":"TESTARE:",
"##showing_agamemnon_aeschylus##":"Uppför: 'Annales', av Tacitus",
"##showing_antigone_sophocles##":"Uppför: Homeros grekiska tragedier",
"##showing_thecrito_plato##":"Uppför: 'Oidipus', av Sofokles",
"##showing_lisistrata_aristopanes##":"Uppför: 'Vergilius dikter'",
"##showing_odyssey_homer##":"Uppför: 'Platons filosofi'",
"##shipyard_info##":"Med några vagnslaster timmer och tillräckligt med arbetare bygger fartygsvarvet fiskebåtar till stadens fiskehamnar.",
"##patrician_average_life##":"Här i min bekväma villa anser jag livet i staden vara mycket bra.",
"##current_game_speed_is##":"Nuvarande spelhastighet",
"##increase_trading_title##":"Begär ändringar",
"##a_price_rise_title##":"Prisändringar",
"##mainmenu_plname##":"Ändra namn
",
"##adjust_exact##":"Ställ in den exakta summa du vill donera",
"##adjust_tax_rate##":"Justera skattenivån i staden",
"##wharf_full_work##":"Med fullt antal anställda lassar och lossar vi med maximal hastighet.",
"##dock_full_work##":"Vi har full arbetsstyrka och kommer att kunna lasta och lossa inkommande fartyg.",
"##wt_immigrant##":"Immigrant",
"##emperor_favour_20##":"Kejsaren är så otroligt nöjd att han talar om att utnämna dig till sin arvinge.",
"##city_still_in_debt_text##":"Kjesaren är rasande på dig för att du fortfarande är skylldig Rom pengar. Han ger dig 12 månader till att betala skulden. Annars kommer du straffas ordentligt.",
"##emperor_favour_18##":"Kejsaren är utom sig av glädje över vad du gjort.",
"##emperor_favour_17##":"Kejsaren är extremt entusiastisk över vad du gjort.",
"##emperor_favour_00##":"Kejsaren är rasande på dig.",
"##emperor_favour_12##":"Kejsaren är tillfreds med dig.",
"##emperor_favour_14##":"Kejsaren är mycket entusiastisk över vad du gjort.",
"##emperor_favour_05##":"Kejsaren är extremt missnöjd med dig.",
"##emperor_favour_02##":"Kejsaren är vansinnigt arg på dig.",
"##emperor_favour_07##":"Kejsaren är missnöjd med dig.",
"##emperor_favour_09##":"Kejsaren är tveksam vad gäller dig.",
"##emperor_favour_08##":"Kejsaren är något missnöjd med dig.",
"##emperor_limit_houseupgrade##":"Kejsaren har begränsat uppgraderingar av husen i denna stad",
"##emperor_favour_13##":"Kejsaren är mycket nöjd med vad du gjort.",
"##emperor_favour_06##":"Kejsaren är mycket missnöjd med dig.",
"##emperor_favour_03##":"Kejsaren är mycket arg på dig.",
"##emperor_favour_16##":"Kejsaren är entusiastisk över vad du gjort.",
"##emperor_favour_11##":"Kejsaren tror du kan bevisa dig värdefull .",
"##emperor_favour_04##":"Kejsaren är arg på dig.",
"##emperor_favour_15##":"Kejsaren är nöjd med vad du gjort.",
"##emperor_favour_01##":"Kejsaren är så otroligt arg att han talar om att landsförvisa dig.",
"##emperor_favour_19##":"Kejsaren är mer än tillfreds med vad du gjort.",
"##imperial_reminder##":"Kjeserlig påminnelse",
"##emperor_request_money##":"Kjesare efterfrågar pengar",
"##emperor_request##":"Kjesare efterfrågar varor",
"##emperor##":"Imperiet",
"##import_fn##":"Importer",
"##import##":"Importerar",
"##trade_btn_import_text##":"Importerar",
"##city_zoominv_on##":"Inverterad zoom: På",
"##city_zoominv_off##":"Inverterad zoom: Av",
"##adve_industry_and_trade##":"Industri och handel",
"##engineer##":"Ingenjör",
"##wt_engineer##":"Ingenjör",
"##adve_engineers##":"Konstruktion",
"##extm_engineering_tlp##":"Ingenjörsbyggnader",
"##engineering_post##":"Ingenjörspostering",
"##engineering_post_info##":"Ingenjörer är mycket respekterade yrkesmän, och det är alltid stor efterfrågan på deras tjänster. Konstant underhåll förhindrar att byggnaderna faller samman.",
"##ready_to_game##":"Redo att spela",
"##hippodrome##":"Hippodrom",
"##ovrm_hippodrome##":"Hippodrom",
"##hippodromes##":"Hippodromer",
"##use_and_trade_resource##":"Använder och byteshandlar med denna vara",
"##citychart_population##":"Historia",
"##caesarea_win_text##":"Så Caesareas förre ståthållare ska alltså få behålla livet? Att rädda staden ur krisen är verkligen en bedrift. Jag kanske ska låta dig välja vilket land vi ska utvisa honom till.",
"##this_year##":"Så här långt detta året",
"##wn_judaean##":"Judeér",
"##judaean_warrior##":"En judéisk soldat",
"##etertadv_as_city_grow_you_need_more_entert##":"Medborgare som söker tidsfördriv har allt vad de behöver. Men i takt med att staden växer måste du förse dem med mer storslagen form av underhållning.",
"##month_7_short##":"Juli",
"##month_6_short##":"Juni",
"##to_trade_advisor##":"Till handelsrådgivaren",
"##walls_need_a_gatehouse##":"Murar behöver grindstugor, så att vandringsmän och handelsmän kan komma och gå som de vill.",
"##barracks##":"Förläggningar",
"##mainmenu_dlc_main##":"Hur man bygger Rom",
"##romeGuard_so_hungry##":"Hur ska en soldat kunna slåss utan mat?",
"##miletus_win_text##":"Precis som jag förväntade mig har exemplet Miletus redan inspirerat andra östliga städer att inleda förhandlingar om att ingå i imperiet. Din erfarenhet av fisket har blivit en läxa för alla mina ståthållare!",
"##patrician_high_workless##":"Detta är skandalöst. Jag har aldrig sett så många arbetslösa plebejer.",
"##capua_title##":"Capoue: une province pacifique",
"##extm_empire_tlp##":"Global karta",
"##empire_map##":"Gå till imperiet",
"##carthago_title##":"Carthago: une province dangereuse",
"##carthaginian_soldier##":"En karthagisk soldat",
"##wn_carthaginians##":"Karthager",
"##earthquake_text##":"Katastrof! Till och med gudarna är chockade. En jordbävning som sväljer allt i sin väg. Hoppas det går bra, reparera alla skador när det slutar.",
"##quaestor##":"Kvestor",
"##wn_celts##":"Kelter",
"##caesarea_title##":"Césarée: province équitablement pacifique",
"##wrath_of_mercury_description##":"Mercury kokar av ilska. Brinnande stenar faller från himlen, som förstör byggnader och dess innehåll!",
"##city_cyrene##":"Cyrene",
"##clerk##":"Bokhållare",
"##clinic##":"Klinik",
"##ovrm_doctor##":"Klinik",
"##clinics##":"Kliniker",
"##londinium_win_text##":"Vid Jupiter! Vildarna i Britannia har aldrig sett Londiniums like. Claudius, som visade öborna de romerska svärdens vassa eggar för många år sedan, ler säkert mot oss från sin himmel.",
"##smcurse2_of_venus_description##":"När Venus är missnöjd sänker hon medborgarnas sinnesstämning. En del säger att hon för med sig sjukdomar.",
"##military_academy_patrly_workers##":"När nya soldater har avslutat sin utbildning i förläggningen kommer de hit för att förbättra och finslipa sina färdigheter. Det går dock först när vi har fått tillräckligt med personal.",
"##middle_fest_description##":"När 1 dagsfesten närmar sig sitt slut, börjar invånare återvända hemåt, trötta men glada. Medan din valda gud ler åt dem alla.",
"##colloseums##":"Colosseum",
"##colloseum##":"Colosseum",
"##colloseum_info##":"Colosseum och amfiteatrar behöver alltid nya gladiatorer för att ersätta förlorarna.",
"##ovrm_colloseum##":"Colleseum",
"##well##":"Brunn",
"##column_info##":"Kolonnformation",
"##ovrm_commerce##":"Handel",
"##consul##":"Konsul",
"##mainmenu_dlc_concepts##":"Begrepp",
"##spear##":"Spjut",
"##fort_javelin##":"Kastspjut",
"##high_bridge##":"Fartygsbro",
"##corinthus##":"Corinthus",
"##extreme_fire_risk##":"Extrem brandrisk",
"##sldr_extremely_scared##":"Extremt rädd",
"##sldh_health_strongest##":"Extremt stark",
"##extm_mission_tlp##":"Titel på provinskarta.",
"##fortification##":"Befästning",
"##blood_sports_add_spice_to_life##":"Blodsporter ger krydda åt alla.",
"##lgn_rabbits##":"Kaninerna",
"##gladiator_pit_bad_work##":"Jag har ingen personal utöver mig själv. Jag kan inte arbeta under dessa förhållanden! Som bäst kan jag utbilda en gladiator var tredje månad.",
"##lion_pit_bad_work##":"Jag har ingen personal utöver mig själv. Jag kan inte arbeta under dessa förhållanden! Som bäst kan jag leverera ett lejon på tre månader.",
"##actorColony_bad_work##":"Jag har ingen personal utöver mig själv. Jag kan inte arbeta under dessa förhållanden! Som bäst kan jag utbilda en skådespelare på tre månader.",
"##chatioteer_school_bad_work##":"Jag har ingen personal utöver mig själv. Jag kan inte arbeta under dessa förhållanden! Jag kan bara bygga en vagn på tre månader.",
"##cartPusher_need_workers##":"Vart man än kommer i staden finns det lediga arbeten.",
"##senatepp_clt_rating##":"Kultur",
"##wndrt_culture##":"Kultur",
"##emw_bought##":"Köpt",
"##romechastener_attack_title##":"Legioner anfaller",
"##emperror_legion_at_out_gates##":"En legion av kejsarens trupper står vid portarna",
"##wt_legioanry##":"Legionär",
"##lumber_mill##":"Brädgård",
"##years##":"Sädesmagasin lagrar",
"##lindum_title##":"Lindum: en extremt farlig provins",
"##line_formation_title##":"Linjeformation",
"##prefecture_full_work##":"För närvarande är vår tjänstgöringslista full. Våra prefekter är alltid ute och patrullerar gatorna.",
"##governor_salary_title##":"Personlig inkomst",
"##pn_salary##":"Personlig inkomst",
"##no_room_for_citizens##":"för många",
"##wharf_info##":"Båtar avseglar från fartygsvarvet och hämtar sina besättningar här. Varje fiskehamn kan betjäna en fiskebåt.",
"##londinium_title##":"Londinium: une province pacifique",
"##meadow_caption##":"Äng",
"##lugdunum_title##":"Lugdunum: une province pacifique",
"##lutetia_title##":"Lutetia: une province dangereuse",
"##road_paved_title##":"En finare typ av väg",
"##animal_contests_run##":"Djurtävlingarna pågår ytterligare",
"##colloseum_haveno_animal_bouts##":"Inga djurkamper för närvarande",
"##lionNusery##":"Lejonhus",
"##lgn_lions##":"Lejonen.",
"##venus_desc##":"Kärlek",
"##dock_no_workers##":"Vi har inga hamnarbetare och kan därför inte lasta eller lossa några fartyg som kommer till hamnen.",
"##bathlady_so_hungry##":"Folk har inte ätit på så länge att deras revben börjar sticka ut, vilket syns på badhuset.",
"##more_4_month_from_festival##":"Människor talar fortfarande varmt om din senaste festival.",
"##citizens_grumble_lack_festivals_held##":"Medborgarna klagar över bristen på festivaler i din stad.",
"##doctor_so_hungry##":"Folk är undernärda, men det saknas mat att bota det med.",
"##more_16_month_from_festival##":"Människorna kommer inte längre ihåg den sista festivalen som hölls i staden.",
"##more_31_month_from_festival##":"Människorna kommer inte längre ihåg den sista festivalen som hölls i staden.",
"##people_leave_city_some##":"Människor lämnar staden",
"##people_leave_city_low_wage##":"Människor beger sig av på jakt efter högre löner",
"##people_leave_city_insane_tax##":"Människor lämnar staden på grund av dina höga skatter",
"##road_paved_text##":"Människor föredrar torg!",
"##migration_peoples_arrived_in_city##":"Människor immigrerar till staden",
"##we_produce_less_than_eat##":"Dina invånare äter mer mat än de producerar",
"##month_5_short##":"Maj",
"##macedonian_soldier##":"En makedonisk soldat",
"##small_villa##":"Liten villa",
"##small_shack##":"Liten koja",
"##small_tent##":"Litet tält",
"##status_small##":"Liten staty",
"##small_hovel##":"Litet skjul",
"##small_hut##":"Litet hus",
"##school_info##":"Barn måste gå i stadsdelsskolorna för att lära sig grunderna i läsning, skrivning och retorik om de skall kunna växa upp till produktiva vuxna.",
"##small_temples##":"Små tempel",
"##bldm_temple##":"Små tempel",
"##small_palace##":"Litet palats",
"##small_domus##":"Liten Insulae",
"##small_festival##":"Liten festival",
"##small##":"Litet",
"##delivery_boy##":"Springpojke",
"##month_3_short##":"Mar",
"##army_marker##":"Armémarkör",
"##god_mars_short##":"Mars",
"##wrath_of_mars_text##":"Mars börjar bli arg på dig. Le om du vågar. Fastän du inte har några millitärastyrkor idag. Mars blir inte så lätt förolämpad. Va vaksam!
",
"##smallcurse_of_mars_failed_text##":"Mars är vrede med dig. Skratta om du inte är rädd, eftersom även idag kan du inte föra krig, kommer Mars inte glömma förolämpningar tillfogat honom. Akta dig!",
"##smallcurse_of_mars_title##":"Mars är upprörd",
"##smallcurse_of_mars_text##":"Mars vakar över soldater och belönar tapperhet i fält. Ingen man vågar kämpa utan Mars välsignelse.",
"##smallcurse_of_mars_text##":"Mars, soldaternas beskyddare och segerförlänare, är missnöjd. Dina soldater fruktar att de kommer att förlora ett stort slag om han inte blidkas.",
"##oil##":"Olja",
"##oil_factory_stock##":"Olja",
"##oil_workshop##":"Oljepresseri",
"##massilia_title##":"Massilia: une province pacifique",
"##chatioteer_school_info##":"De hantverkare som arbetar här bygger snabba, kraftiga vagnar och utbildar förarna. Kapplöpningarna i hippodromen är mycket populära.",
"##cartpusher_cant_unload_goods_in_factory##":"...ta emot dem. Jag har hört att de behöver mer arbetskraft.",
"##bldm_factory##":"Verkstäder",
"##furniture##":"Möbler",
"##furniture_workshop##":"Möbelsnickeri",
"##mediolanum_title##":"Mediolanum: province très dangereux",
"##balance_between_migration##":"Det är lika många som kommer till, respektive lämnar staden",
"##gmenu_file##":"Arkiv",
"##emigrant_thrown_from_house##":"Jag har blivit utkastad från mitt hem!",
"##mercury##":"Mercury",
"##smcurse_of_mercury_title##":"Merkurius är upprörd",
"##smallcurse_of_mercury_failed_title##":"Mercury is upprörd",
"##smallcurse_of_mercury_title##":"Mercury is upprörd",
"##smallcurse_of_mercury_description##":"Merkurius, gudarnas budbärare och handelsmännens beskyddare, är missnöjd. Dina handelsmän fruktar att hans beskydd viker.",
"##native_center_info##":"Mötesplats för lokalbefolkningen",
"##unhandled_key_value_19##":"Plats för en nyligen inträffad sammandrabbning med invaderande barbarer",
"##month##":"Mes",
"##month_to_comply##":"Mes",
"##months##":"Människor",
"##rqst_month_2_comply##":"Människor",
"##months_to_comply##":"Människor",
"##months_until_victory##":"Månader till seger",
"##months_until_defeat##":"Månader till nederlag",
"##wt_romeSpearman##":"Spjutkastare",
"##miletus_title##":"Milet: province largement pacifique",
"##warning_hippodrome_access##":"Detta hus har inte passerats av en körsven på ett tag. Det kommer snart att förlora tillgång till hippodrom",
"##warning_amphitheater_access##":"Detta hus har inte passerats av en gladiator på ett tag. Det kommer snart att förlora tillgång till amfiteater",
"##warning_colloseum_access##":"Detta hus har inte passerats av en lejontämjare på ett tag. Det kommer snart att förlora tillgång till colosseum",
"##avesome_amphitheater_access##":"Detta hus passerades nyligen av en gladiator. Det kommer att ha tillgång till amfiteater under lång tid framåt",
"##avesome_theater_access##":"Detta hus passerades nyligen av en skådespelare. Det kommer att ha tillgång till teater under lång tid framåt",
"##avesome_library_access##":"Detta hus har nyligen passerats av en bibliotekarie. Det kommer att ha tillgång till bibliotek under lång tid framåt",
"##avesome_hippodrome_access##":"Detta hus har nyligen passerats av en körsven. Det kommer att ha tillgång till hippodrom under lång tid framåt",
"##avesome_clinic_access##":"Detta hus passerades nyligen av en läkare. Det kommer att ha tillgång till en klinik under lång tid framåt",
"##awesome_barber_access##":"Detta hus passerades nyligen av en barberare. Det kommer att ha tillgång till en barberare under lång tid framåt",
"##avesome_colloseum_access##":"Detta hus passerades nyligen av en lejontämjare. Det kommer att ha tillgång till ett colosseum under lång tid framåt",
"##avesome_college_access##":"Detta hus passerades nyligen av en lärare. Det kommer att ha tillgång till högskola under lång tid framåt",
"##avesome_hospital_access##":"Detta hus passerades nyligen av en kirurg. Det kommer att ha tillgång till sjukhus under lång tid framåt",
"##avesome_school_access##":"Detta hus passerades nyligen av ett skolbarn. Det kommer att ha tillgång till skola under lång tid framåt",
"##awesome_baths_access##":"Detta hus passerades nyligen av en badhusarbetare. Det kommer att ha tillgång till badhus under lång tid framöver",
"##senatepp_peace_rating##":"Fred",
"##wt_missionary##":"Missionär",
"##missionaryPost##":"Inhemsk mission",
"##taxCollector_high_workless##":"Jag ogillar det här stället. Arbetslösheten är för hög.",
"##emigrant_no_work_for_me##":"Jag har fått nog av detta ställe. Det finns inget arbete här.",
"##emigrant_no_home##":"Jag har ingenstans att bo.",
"##taxСollector_much_tax##":"Jag älskar att driva in skatt från rika hus som dessa.",
"##legionary_low_salary##":"Jag får inte tillräckligt bra betalt för att slåss!",
"##healthadv_some_regions_need_barbers##":"Fler områden i staden kräver nu barberare. I takt med att din stad blir allt mer välbeställd kommer fler att ha tid till rakning och klippning!",
"##much_plebs##":"Den höga koncentrationen av boende i slumområden i din stad gör att den ser fattig ut.",
"##max_available##":"Underhåller",
"##centurion_send_army_to_player##":"Mitt tålamod är slut. Då du fortfarande inte har bra relation med Kjesaren, måste jag tyvärr utföra mina order, oavsett hur otäcka de är. Ge upp nu eller bered dig på konsikvenserna!",
"##freespace_for##":"Utrymme för",
"##my_rome##":"Mitt Rom",
"##pestilence_event_title##":"Farsot",
"##neptune_desc##":"Havet",
"##neptune_despleasure_tip##":"Sjömän finner att Neptunus är en ombytlig gud även om han blidkas. Väck inte Neptunus vrede, om du önskar bedriva handel över vattnet.",
"##bridge##":"Bro",
"##bridges##":"Broar",
"##road_paved_caption##":"Stenbelagdväg",
"##plaza_caption##":"Torg",
"##plaza##":"Torg",
"##marble##":"Marmor",
"##quarry##":"Marmorbrott",
"##gmsndwnd_theme_sound##":"Musik",
"##mainmenu_dlc_soundtrack##":"Teman",
"##music##":"MUSIK:",
"##floatsam_enabled##":"Vrakgods på?",
"##priest_gods_angry##":"Vi är i fara! Staden visar ingen respekt för gudarna.",
"##wait_for_fishing_boat##":"Vi vänta för närvarande på att ett varv skall bygga oss en fiskebåt.",
"##prefecture_bad_work##":"Vi arbetar endast med kontorspersonal. Det går ofta en hel månad utan att vi sänder en prefekt ut på gatorna.",
"##missionaryPost_full_work##":"Vi arbetar på att civilisera lokalbefolkningen. Genom att lära dem grunderna i latin hoppas vi uppmuntra dem att arbeta med oss, istället för emot oss.",
"##barracks_no_weapons##":"Vi kan utbilda stödtrupper mycket snabbt, men utan vapenupplag kan vi inte utbilda några nya legionärer.",
"##dock_busy_patrly_workers##":"Vi betjänar det förtöjda fartyget, trots att vi inte har tillräckligt med anställda, så det kommer att ta längre tid än det borde.",
"##dock_busy_bad_work##":"Vi betjänar det förtöjda fartyget, men har för få hamnarbetare, detta kommer att ta tid.",
"##barracks_full_work##":"Vi utbildar nya soldater med maximal effektivitet och vi har vapen för att utbilda alla typer av soldater.",
"##barracks_need_some_workers##":"Pga. personalbrist utbildar vi nya soldater långsammare än vanligt men vi har de vapen som krävs för att utbilda alla typer av soldater.",
"##getting_reports_about_enemies##":"Vi får rapporter om fiender som närmar sig staden",
"##restocking_fishing_boat##":"Vi förbereder för närvarande vår fiskebåt för att segla ut igen. Hur snabbt det går beror på hur många anställda vi har.",
"##we_eat_more_thie_produce##":"Vi äter mer än vi producerar",
"##we_eat_much_then_produce##":"Vi äter mycket mer än vi producerar",
"##we_eat_some_then_produce##":"Vi äter något mer än vi producerar",
"##we_produce_some_than_eat##":"Vi producerar lagom för att livnära alla",
"##we_produce_much_than_eat##":"Vi producerar mycket mer än vi äter",
"##we_produce_more_than_eat##":"Vi producerar något mer än vi äter",
"##engineering_post_bad_work##":"Vi arbetar med minimistyrka. Vi kan knappt sända ut en ingenjör per månad på fältet.",
"##lion_pit_work##":"Det är med nöje vi tillkännager att vi, med full sysselsättning, kan leverera upp till fyra nya lejon varje månad.",
"##actorColony_full_work##":"Det är med nöje vi tillkännager att vi, med full sysselsättning, kan hjälpa upp till fyra nya skådespelare varje månad.",
"##charioteer_school_full_work##":"Det är med nöje vi tillkännager att vi, med full sysselsättning, kan slutföra upp till fyra nya vagnar varje månad.",
"##gladiator_pit_full_work##":"Det är med nöje vi tillkännager att vi, med full sysselsättning, utbildar upp till fyra nya gladiatorer varje månad.",
"##enemies_very_easy##":"Vi ska nog skrämma bort veklingarna snabbt.",
"##enemies_very_hard##":"Vi ska göra vårt bästa, men även romerska soldater får svårt att besegra den här fienden.",
"##lionTamer_low_entertainment##":"Leo och jag slåss dygnet runt och ändå har folk tråkigt. Det finns helt enkelt inte tillräckligt med artister här.",
"##build_fishing_boat##":"Vi bygger båtar på beställning från en fiskehamn i staden.",
"##militaryAcademy_full_work##":"Vi förser nya rekryter från stadens förläggningar med den ytterligare utbildning de kräver för att fungera bra i en modern romersk armé.",
"##meat##":"Kött",
"##ad##":"eKr",
"##age_ad##":"eKr",
"##need_trainee_charioteer##":"Det finns inga kapplöpningsvagnar i din hippodrom. Anskaffning av sådana skulle avsevärt förbättra villkoren för befolkningen, som ivrigt söker mer underhållning.",
"##no_goods_for_request##":"Du har inte tillräckligt med varor i dina handelsmagasin",
"##scholar_gods_angry##":"Hjälp! Gudarna är vreda. De kommer att straffa oss.",
"##marketLady_no_food_on_market##":"Marknaden har slut på livsmedel, så jag är på väg hem.",
"##wine_workshop_full_work##":"Denna vingård har alla anställda den behöver och arbetar fullt ut med att producera vin.",
"##wine_workshops_need_some_workers##":"Denna vingård är underbemannad och det tar mycket längre tid att producera vin än vad det borde.",
"##wine_workshop_no_workers##":"Denna vingård har inga anställda. Produktionen har upphört.",
"##wine_workshop_slow_work##":"Mycket få människor arbetar vid denna vingård. Som resultat är vinproduktionen långsam.",
"##clear_land_text##":"Detta landområde kan byggas på efter behov. Det ger fri passage både åt egna soldater och åt fiendesoldater.",
"##lumber_mill_full_work##":"Denna brädgård har alla anställda den behöver. Den arbetar fullt ut med att såga timmer.",
"##lumber_mill_patrly_workers##":"Denna brädgård är underbemannad, och det tar längre tid att såga virke än vad det borde.",
"##lumber_mill_no_workers##":"Denna brädgård har inga anställda. Produktionen har upphört.",
"##lumber_mill_slow_work##":"Mycket få människor arbetar vid den här brädgården. Som resultat är timmerproduktionen långsam.",
"##oil_workshop_slow_work##":"Mycket få människor arbetar vid denna olivpress. Som resultat är oljeproduktionen långsam.",
"##fig_farm_full_work##":"Denna fruktträdgård har alla anställda den behöver. Träden dignar av mogen frukt.",
"##olive_farm_full_work##":"Denna lund har alla anställda den behöver. Trädgrenarna dignar med tunga lass av oliver.",
"##meat_farm_full_work##":"Denna farm har alla anställda den behöver, och dess djurstam är fet och stor.",
"##vegetable_farm_need_some_workers##":"Denna lantgård är underbemannad. Vissa av dess grönsaker kommer att ruttna på åkern.",
"##olive_farm_patrly_workers##":"Denna lund är underbemannad. Det tar längre tid att plocka oliverna än vad det borde.",
"##wheat_farm_need_some_workers##":"Denna lantgård är underbemannad. Arbetarna kan inte så alla de fält som finns.",
"##meat_farm_need_some_workers##":"Denna farm är underbemannad. Svinen har små kullar, som växer långsamt.",
"##fig_farm_need_some_workers##":"Denna fruktträdgård är underbemannad. Den producerar mindre frukt än vad den borde.",
"##meat_farm_no_workers##":"Denna farm har inga anställda, och alla djuren har flytt eller dött.",
"##olive_farm_no_workers##":"Denna lantgård har inga anställda. Inget har planterats.",
"##vegetable_farm_no_workers##":"Denna lantgård har inga anställda. Inget har planterats.",
"##wheat_farm_no_workers##":"Denna lantgård har inga anställda. Jorden ligger i träda.",
"##fig_farm_no_workers##":"Denna fruktträdgård har inga anställda. Produktionen har upphört.",
"##unhandled_key_value_17##":"Denna lund har inga anställda. Produktionen har upphört.",
"##meat_farm_slow_work##":"Mycket få människor arbetar på den här farmen. Som resultat är köttproduktionen långsam.",
"##vegetable_farm_full_work##":"Denna lantgård har alla anställda det behöver. Grönsaker växer här i överflöd.",
"##wheat_farm_full_work##":"Denna lantgård har alla anställda det behöver. Den får maximum avkastning på sin areal.",
"##vinard_full_work##":"Denna odling har alla anställda den behöver. Vinrankorna är tunga med stora, saftiga druvor.",
"##vinard_need_some_workers##":"Denna odling är underbemannad. Det tar längre tid att producera druvor än vad det borde.",
"##vinard_no_workers##":"Denna odling har inga anställda. Produktionen har upphört.",
"##vinard_slow_work##":"Mycket få människor arbetar på denna odling. Som resultat är druvproduktionen långsam.",
"##trouble_hippodrome_no_charioters##":"Denna hippodrom kör inga kapplöpningar. Den behöver körsvenner.",
"##trouble_hippodrome_full_work##":"Denna hippodrom har ofta spännande kapplöpningar, som ger mycket nöje åt lokalbefolkningen.",
"##clay_pit_full_work##":"Detta lertag har alla anställda det behöver, och arbetar fullt ut med att producera lera.",
"##quarry_full_work##":"Detta brott har alla anställda det behöver, det arbetar fullt ut med att producera marmor.",
"##clay_pit_patrly_workers##":"Detta lertag är underbemannat, och det tar längre tid att producera leran än vad det borde.",
"##quarry_patrly_workers##":"Detta brott är underbemannat, och det tar längre tid än det borde att producera marmorn.",
"##clay_pit_no_workers##":"Detta lertag har inga anställda. Produktionen har upphört.",
"##quarry_no_workers##":"Detta brott har inga anställda. Produktionen har upphört.",
"##quarry_slow_work##":"Mycket få människor arbetar vid detta lertag. Som resultat är lerproduktionen långsam.",
"##quarry_patrly_workers##":"Mycket få människor arbetar vid det här brottet. Som resultat är marmorproduktionen långsam.",
"##oil_workshop_full_work##":"Denna olivpress är fullt bemannad och producerar rikliga mängder olja av hög kvalitet.",
"##oil_workshop_need_some_workers##":"Denna olivpress behöver fler arbetare för att nå sin fulla potential för oljeproduktion.",
"##oil_workshop_no_workers##":"Denna olivpress har inga anställda och kommer inte att producera olja.",
"##iron_mine_full_work##":"Detta brott har alla anställda det behöver, och arbetar fullt ut med att producera järn.",
"##iron_mine_patrly_workers##":"Detta brott är underbemannat. Det tar längre tid än normalt att producera järnet.",
"##iron_mine_no_workers##":"Detta brott har inga anställda. Produktionen har upphört.",
"##iron_mine_slow_work##":"Mycket få människor arbetar vid det här brottet. Som resultat är järnproduktionen långsam.",
"##market_search_food_source##":"Denna marknad har köpmän men de söker för närvarande efter en källa till livsmedel som kan säljas.",
"##water_srvc_fountain_and_well##":"Detta område har tillgång till en reservoar via rörledning och dricksvatten från en brunn eller fontän",
"##teacher_high_workless##":"Bara jag inte förlorar jobbet. Arbetslösheten är så hög att jag inte skulle få ett nytt.",
"##fort_horse##":"Stödtrupp - Ridande",
"##press_escape_to_exit##":"Högerklicka för att avsluta",
"##restart_mission_tip##":"Klicka här för att återuppbygga denna provins",
"##set_mayor_salary##":"Klicka här för att fastställa din personliga lön",
"##click_here_that_use_it##":"Klicka här för att stänga av hamstring",
"##legion_formation_tooltip##":"Klicka här för att ändra legionens formation",
"##click_here_that_stacking##":"Klicka här för att hamstra",
"##request_btn_tooltip##":"Klicka här för att sända iväg begäran",
"##give_money_tip##":"Klicka här för att donera pengar till staden",
"##go_to_problem##":"Klicka här för att gå till detta problemområde",
"##click_here_to_talk_person##":"Klicka här för att tala med denna person",
"##advice_at_culture##":"Klicka här för information om din kulturställning",
"##wndrt_favor_tooltip##":"Klicka här för information om din popularitetsställning",
"##wndrt_peace_tooltip##":"Klicka här för information om din fredsställning",
"##wndrt_prosperity_tooltip##":"Klicka här för information om din välståndsställning",
"##empbutton_tooltip##":"Klicka här för att fastställa en prioritet för denna arbetskraftskategori",
"##land_route##":"Landväg",
"##having_some_slums_lack_migration##":"Att ha slumområden förhindrar immigration",
"##taxes##":"Inkasserade skatter",
"##ovrm_tax##":"Skatter",
"##engineering_post_slow_work##":"Vi är kraftigt underbemannade och har en tidslucka på två veckor mellan ingenjörernas rundor.",
"##forum_1_slow_work##":"Vi är kraftigt underbemannade och har en lucka på två veckor innan indrivarna ger sig ut.",
"##chatioteer_school_slow_work##":"Vi lider av svår personalbrist, och kommer att få kämpa för att bygga en enda ny vagn under de kommande två månaderna.",
"##actorColony_slow_work##":"Vi lider av svår personalbrist, och kommer att få kämpa för att utbilda en ny skådespelare under de kommande två månaderna.",
"##prefecture_patrly_workers##":"Vi är underbemannade, och har farliga luckor på upp till en vecka i vår tjänstgöringslista.",
"##barracks_bad_weapons_slow_workers##":"Vi är underbemannade och saknar vapen, vi kan bara långsamt utbilda stödtrupper.",
"##engineering_post_patrly_workers##":"Vi har för lite personal, så vi måste vänta en vecka innan våra ingenjörer är tillbaka i tjänst.",
"##actorColony_need_some_workers##":"Vi är något underbemannade, och kan därför endast utbilda två nya skådespelare per månad.",
"##lion_pit_need_some_workers##":"Vi är något underbemannade, och kan därför endast leverera två nya lejon i månaden.",
"##gladiator_pit_need_some_workers##":"Vi är något underbemannade, och kan därför endast utbilda två nya gladiatorer i månaden.",
"##charioteer_school_need_some_workers##":"Vi är något underbemannade, och kan därför endast tillverka två nya vagnar per månad.",
"##barracks_bad_weapons_need_some_workers##":"Vi saknar några anställda och utbildar soldater långsammare än vanligt. Utan vapenupplag kan vi inte utbilda några nya legionärer.",
"##prefecture_need_some_workers##":"Vi har lite ont om prefekter. Vi har luckor på en dag eller två i vår täckning.",
"##gladiator_pit_slow_work##":"Vi lider av svår personalbrist, och kommer att få kämpa för att utbilda en ny gladiator under de kommande två månaderna.",
"##lion_pit_slow_work##":"Vi lider av svår personalbrist, och kommer att få kämpa för att leverera ett enda lejon under de kommande två månaderna.",
"##heading_to_city_warehouses##":"På väg mot stadens handelsmagasin",
"##people##":"denarer",
"##peoples##":"denarer",
"##pop##":"Inv",
"##advlegion_norequest##":"Vi har inte fått någon begäran om hjälp från imperiet",
"##mission_wnd_population##":"Befolkning",
"##population##":"Befolkning",
"##winning_population##":"Vinnande befolkning",
"##advpopulation_title_census##":"Befolkning - Folkräkning",
"##advpopulation_title_society##":"Befolkning - Samhälle",
"##advpopulation_title_population##":"Befolkning - Historia",
"##lowgrade_housing_want_better_conditions##":"Invånarna i dåliga bostäder vill ha bättre villkor",
"##population_registered_as_taxpayers##":"av befolkningen är skatteskrivna",
"##advchief_sentiment##":"Stämning",
"##gmenu_options##":"Alternativ",
"##mainmenu_options##":"Alternativ",
"##options##":"Inställning",
"##city_options##":"Stadalternativ",
"##mainmenu_sound##":"Ljudinställningar",
"##sound_settings##":"Ljudinställningar",
"##game_sound_options##":"Ljudalternativ",
"##city_settings##":"Stadinställningar",
"##speed_settings##":"Hastighetsinställningar",
"##game_speed_options##":"Hastighetsinställningar",
"##mainmenu_video##":"Bildskärmsinställningar",
"##screen_settings##":"Bildskärmsinställningar",
"##start_condition##":"Startvillkor",
"##replay_game##":"Börja om denna karta",
"##start_this_map##":"Starta denna karta",
"##mainmenu_startcareer##":"Ny karriär",
"##devastate_warehouse##":"BÖRJA tömma magasin",
"##empiremap_our_city##":"Vår stad!",
"##engineering_post_ready_for_work##":"Vår ingenjör förbereder sig för att ge sig av.",
"##engineering_post_on_patrol##":"Vår ingenjör är ute och arbetar.",
"##out_legion_back_to_city##":"Vår legion marscherar tillbaka till vår stad",
"##out_legion_go_to_location##":"Vår legion marscherar för att rädda en av rikets städer",
"##prefecture_ready_for_work##":"Vår prefekt förbereder sig för sin tjänst.",
"##prefecture_on_patrol##":"Vår prefekt är ute och patrullerar.",
"##forum_1_ready_for_work##":"Vår indrivare förbereder sig för att ge sig av.",
"##forum_1_on_patrol##":"Vår indrivare är ute på inspektion.",
"##wharf_our_boat_fishing##":"Vår fiskebåt befinner sig vid fiskevattnet och fångar just nu fisk.",
"##wharf_our_boat_return##":"Vår båt seglar mot hamn.",
"##wharf_out_boat_ready_fishing##":"Vår fiskebåt seglar ut till fiskevattnen.",
"##wharf_out_boat_return_with_fish##":"Vår fiskebåt seglar tillbaka från fiskevattnen med sin fångst.",
"##dock_cart_returning_from":"Vår vagn återvänder från en leverans.",
"##dock_cart_taking_goods##":"Vår vagn för varorna till annan plats.",
"##dock_cart_wait##":"Vår vagn är här och väntar på nya order.",
"##unhandled_key_value_16##":"Våra trupper behövs på annan plats",
"##unhandled_key_value_15##":"Vi har trupper på annan plats",
"##our_enemies_near_city##":"Våra fiender är inom synhåll från staden",
"##our_foods_level_are_low##":"Våra livsmedelsförråd är små",
"##unhandled_key_value_14##":"Våra män är redo att slå tillbaka barbarattacker.",
"##no_fishplace_in_city##":"Vår fiskebåt hoppas snart kunna hitta en fiskeplats. Det blir svårt att försörja sig om vi inte hittar fisk...",
"##market_about##":"Våra marknader gör imperiets rika håvor tillgängliga för medborgare med pengar. Varje hem behöver tillgång till en marknad, men ingen vill bo intill en.",
"##not_available##":"Ej tillgänglig... ännu!",
"##landmerchant_noany_trade##":"Jag vet inte varför jag tar den här handelsvägen. De köper ingenting och de har inget de vill sälja till mig.",
"##merchant_wait_for_deal##":"Jag vill gärna göra affärer här. Jag älskar att göra en bra affär.",
"##no_visited_by_taxman##":"Ej fått besök av skatteindrivare. Betalar ej skatt",
"##reject##":"Avvisa varor",
"##donot_organize_festival##":"Organisera ingen festival",
"##abwrk_not_working##":"fungerar inte",
"##warehouse_low_personal_warning##":"Underbemannad. Kan endast sända iväg varor, ej ta emot varor",
"##unable_fullfill_request##":"Kan inte fullgöra begäran",
"##need_build_on_free_area##":"Du måste bygga på barmark",
"##last_riots_bad_for_peace_rating##":"Upploppen som nyligen ägde rum i staden har haft negativ inverkan på din fredsställning!",
"##imperial_request_cance_badly_affected##":"Den kejserliga begäran som du nyligen upphävde har skadat din ställning i Rom.",
"##several_crimes_but_area_secure##":"Flera brott har rapporterats här nyligen, men på det hela taget har prefekterna situationen under kontroll",
"##rioter_in_city_text##":"Vandalism härjar på dina gator. De är missnöjda med hur guvernören ignorerat deras klagan på villkoren.",
"##god_displeased##":"Missnöjda",
"##ceres_badmood_info##":"Ceres missnöje är farligt, eftersom hon skyddar folket från dåliga skördar och hungersnöd.",
"##out_of_credit##":"Kredit saknas!",
"##city_fire_text##":"Dåligt underhåll har gjort att det börjat brinna. Just nu sveper elden genom olika områden i staden.",
"##some_fire_risk##":"Viss brandrisk",
"##little_damage_risk##":"Viss risk att kollapsa",
"##god_indifferent##":"Likgiltiga",
"##some_houses_inadequate_entertainment##":"Vissa medborgare klagar över bristande tillgång till underhållning i sina områden. Du kanske behöver erbjuda ett mer varierat utbud, eller kanske bygga fler skådespelarkolonier till dina teatrar.",
"##religionadv_need_third_religion##":"Vissa medborgare vill ha en tredje religion etablerad nära sitt område. De anser att detta skulle attrahera bättre patricierklasser.",
"##academy_info##":"En del ungdomar som går ut skolorna går vidare och studerar avancerad retorik och historia vid högskolan. Alla kulturella medborgare har en akademisk bakgrund.",
"##have_no_access_school_colege##":"Vissa områden kräver bättre tillgång till skolor och högskolor. Endast vissa hus har tillgång till skolor eller högskolor, och detta hindrar områdenas utveckling.",
"##advchief_some_need_baths##":"Vissa medborgare behöver badhus",
"##religionadv_need_second_religion##":"Medborgarna i vissa områden vill ha tillgång till en annan religion nära hemmet. Bristen på religioner hindrar stadens utveckling i vissa områden.",
"##advchief_some_need_library##":"Vissa medborgare vill ha fler bibliotek",
"##advchief_some_need_academy##":"Vissa medborgare vill ha fler skolor",
"##advchief_some_need_doctors##":"Vissa medborgare behöver läkarkliniker",
"##advchief_some_need_hospital##":"Vissa medborgare behöver sjukhus",
"##advchief_some_need_barber##":"Vissa medborgare behöver barberare",
"##healthadv_some_regions_need_bath_2##":"Vissa områden i staden behöver nu tillgång till badhus. Bristen på dessa sanitära anläggningar begränsar byggnadstillväxten i dessa områden.",
"##have_no_access_to_library##":"Tillgång till bibliotek krävs nu i vissa delar av staden. Dina medborgare har tid att läsa. Nu behöver de tillgång till litteratur.",
"##healthadv_some_regions_need_doctors##":"Vissa delar av staden kräver tillgång till en klinik. Utan någon form av hälsovård kommer dessa hus förmodligen inte att växa.",
"##some_houses_need_library_or_colege_access##":"Vissa områden i staden kräver nu skolor och högskolor. Bristen på utbildningsmöjligheter förhindrar byggandet av bättre bostäder i dessa områden.",
"##some_houses_need_better_library_access##":"Vissa områden i staden vill ha bättre tillgång till bibliotek. Välbärgade medborgare tycker om att läsa men vill inte gå långt för att nå biblioteket.",
"##edadv_need_better_access_school_or_colege##":"Bättre skola eller högskola och tillgång till bibliotek skulle förbättra vissa områden i staden. Man skall inte behöva gå långt för att lära sig något!",
"##healthadv_some_regions_need_bath##":"Vissa delar av staden vill ha fler badhus. Vissa hus har tillgång till bad, men andra har det inte, och detta hindrar deras utveckling.",
"##some_soldiers_need_weapon##":"Vissa soldater måste ha tillgång till vapenförråd",
"##advchief_some_need_education##":"Medborgarna kräver mer utbildning",
"##scribemessages_unread##":"Oläst meddelande. Vänsterklicka på detta meddelande för att läsa det.  Högerklicka på detta meddelande för att radera det",
"##smallcurse_of_neptune##":"Neptunus skyddar sjömän och deras skepp från havets faror. Om du gör honom missnöjd riskerar du dina sjömäns liv.",
"##god_neptune_short##":"Guden Neptune...",
"##smallcurse_of_neptune_title##":"Neptunus är upprörd",
"##god_poor##":"Dålig",
"##unhandled_key_value_13##":"Inga problem rapporteras",
"##no_priority##":"Ingen prioritet",
"##no_fire_risk##":"Ingen brandrisk",
"##none_damage_risk##":"Ingen risk för kollaps",
"##trade_btn_notrade_text##":"Gör ej affärer",
"##unhandled_key_value_12##":"Ingen begäran",
"##migration_lessfood_granary##":"Brist på livsmedel i sädesmagasinen minskar immigrationen",
"##migration_empty_granary##":"Brist på mat förhindrar immigration",
"##migration_people_away##":"Brist på arbete driver bort människor",
"##migration_middle_lack_workless##":"Brist på arbete förhindrar immigration",
"##migration_lack_empty_house##":"Brist på husrum begränsar immigrationen",
"##barber_info##":"Ingen civiliserad man visar sig orakad offentligt! Alla medborgare behöver regelbundet besöka en barberare för att kunna avancera i samhället.",
"##shipyard_notneed_ours_boat##":"Det finns för närvarande inga fiskehamnar som behöver våra båtar.",
"##below_average##":"Under medel",
"##low_wage_broke_migration##":"Låga löner förhindrar immigration",
"##low_wage_midlle_migration##":"Låga löner minskar immigrationen till din stad",
"##low_bridge##":"Låg bro",
"##low_fire_risk##":"Liten brandrisk",
"##low_damage_risk##":"Liten risk att kollapsa",
"##unhandled_key_value_10##":"Inga spår av barbarer.",
"##unhandled_key_value_11##":"Inga spår av fienden.",
"##prefect_high_workless##":"Jag har aldrig sett så många arbetslösa!",
"##freehouse_text_noroad##":"Ingen kommer att skapa sig ett hem här eftersom det ligger för långt från närmaste väg. Om ingen väg byggs snart kommer detta område att återgå till öppet landskap.",
"##barracks_info##":"Ingen kan gå med i en romersk legion utan att först komma hit. Alla nya rekryter kommer hit.",
"##unhandled_key_value_9##":"Ingen vill bo i din stad",
"##no_citizens_desire_live_here##":"Inga medborgare vill bo här",
"##ovrm_simple##":"Ingenting",
"##plname_start_new_game##":"Ny karriär",
"##mainmenu_newgame##":"Nytt spel",
"##new_map##":"Ny karta
",
"##valencia_win_text##":"Hispaniens nya huvudstad är precis vad vi behöver för att knyta den avlägsna provinsen tätare till Rom. Genom att krossa etruskerna så totalt försvinner det sista hotet i väst.",
"##barber_so_hungry##":"En hårklippning får dig att glömma hungern. Och det är många hungriga i den här staden.",
"##newcomer_this_month##":"nykomling anlände denna månad",
"##new_governor##":"Den nya guvernören",
"##new_ruler##":"Une nouvelle règle",
"##newcomers_this_month##":"nykomlingar anlände denna månad",
"##wt_cartPusher##":"Vagndragare",
"##month_11_short##":"Nov",
"##wndrt_need##":"Behövs",
"##advemployer_panel_needworkers##":"behöver",
"##city_need_workers_title##":"Behöver fler arbetare",
"##furniture_need##":"Möbler behövs",
"##carthago_preview_mission##":"Numidiskt kavalleri har plågat områdena söder om Thamugadi i många år. Du kan vara säker på att de kommer att pröva din försvarsförmåga också.",
"##numidian_warrior##":"En numidisk soldat",
"##wn_numidian##":"Numidier",
"##amazing_prosperity_this_city##":"Det fantastiska välståndet i den här staden är det stora samtalsämnet i Rom!",
"##gmenu_about##":"Om",
"##smcurse_of_mercury_description##":"Förfärad över ditt bristande intresse för honom har Merkurius med andlig kraft avlägsnat en del varor från dina sädes- eller handelsmagasin.",
"##greatPalace_info##":"De boende i detta palats befinner sig högst upp i det romerska samhället. De saknar inte något. Bara att lyckas hålla dem nöjda är en storartad insats.",
"##floatsam##":"Vrakgods",
"##mainmenu_dlc_wallpapers##":"Bakgrundsbilder",
"##legion##":"Militär",
"##blessing_of_mercury_description##":"Förtjust över din hängivenhet har Merkurius upptäckt bortglömda produkter i ett av stadens sädesmagasin.",
"##advchief_education##":"Utbildning",
"##education_advisor_title##":"Utbildning",
"##education##":"Utbildning",
"##educationBtnTooltip##":"Utbildning",
"##ovrm_educations##":"Utbildning",
"##egift_educated_slave##":"En utbildad slav",
"##extm_education_tlp##":"Utbildningsbyggnader",
"##collapse_immitent##":"Överhängande risk för kollaps",
"##iron_mine_collapse##":"Malmbrott kollapsar",
"##academy_trained##":"Utbildad på högskola",
"##bad_house_quality##":"Den totala kvaliteten på byggnaderna i din stad inverkar negativt på denna ställning.",
"##extm_water_tlp##":"Byggnader förknippade med vatten",
"##health_advisor##":"Byggnader förknippade med hälsa",
"##vegetable##":"Grönsaker",
"##vegetable_farm_info##":"Grönsaker är en viktig del av den balanserad diet som ditt folk behöver för hälsa och glädje. I sädesmagasinen lagras grönsaker för lokal konsumtion, och i handelsmagasinen förvaras överskottet för export.",
"##vegetable_farm##":"Grönsaksodling",
"##wt_sheep##":"Får",
"##beatyfull_insula##":"Storslagen Insulae",
"##ok##":"OK",
"##fullscreen_off##":"Upplösning",
"##month_10_short##":"Okt",
"##olive##":"Oliver",
"##olive_farm_info##":"Oliver är värdefulla för sin olja. Olivpresserierna ger olja för matlagning, belysning, smörjning och konservering.",
"##olive_farm##":"Olivodling",
"##export_btn_tooltip##":"Fastställ den kvantitet av dessa varor som du önskar behålla innan de exporteras",
"##distribution_center##":"Distributionscentral",
"##devastate_granary##":"Töm sädesmagasin",
"##oracle##":"Orakel",
"##oracles_in_city##":"Orakel i staden",
"##oracles##":"Orakel",
"##original_game##":"URSPRUNGLIGA SPELET:",
"##weapons_workshop##":"Vapensmedja",
"##weapons_workshop_info##":"Vapensmeder förvandlar järn till vapen och rustningar, som du kan handla med och göra vinst eller använda för att utrusta dina egna legioner.",
"##weapon##":"Vapen",
"##wrath_of_ceres_description##":"Förgrummad över din brist av respekt mot Ceres, hon ger ditt folk en gräshopsplåga. Det kommer dröja innan dina grödor kan växa igen.",
"##unhandled_key_value_1##":"Stöttepelaren i den romerska armétaktiken. Ger stora fördelar mot anfallande fiender.",
"##landmerchant_say_about_store_goods##":"Försiktigt! Jag önskar att arbetarna skulle ta det lugnt när de lastar mina djur med de varor jag nyss har köpt.",
"##sdlr_bold##":"Modig",
"##empmap_distant_romecity_tip##":"Avlägsen romersk stad",
"##some_houses_need_amph_for_grow##":"Vissa medborgare klagar över bristande tillgång till fritidsanläggningar. Vissa områden i staden kräver mer varierade underhållningsmöjligheter.",
"##entertainment_need_for_upgrade##":"I delar av staden klagar man över frånvaron av fritidsanläggningar. Byggnation av fler platser för underhållning skulle hjälpa utvecklingen i de fattigare områdena.",
"##healthadv_some_regions_need_barbers_2##":"Vissa välbeställda delar av staden vill ha barberare. En lokal barberare ger bättre status åt området.",
"##setup_traderoute_to_import##":"Fastställ en handelsväg för att importera det",
"##new_trade_route_to##":"Ny handelsväg etablerad.",
"##mainmenu_randommap##":"Öppet spel ",
"##open_formation_title##":"Öppen formation",
"##open_formation_text##":"Öppen ordning ger möjlighet att täcka ett brett område, men ger dem ingen formationsfördel.",
"##maximizeBtnTooltip##":"Visa fönster",
"##open_trade_route##":"Öppna handelsväg",
"##emp_open_trade_route##":"Öppna handelsväg",
"##god_excellent##":"Utmärkt",
"##cancel##":"Avbryt",
"##extm_cancel_tlp##":"Avbryt denna operation",
"##disabled_draw_salary_for_free_reign##":"Senaten förbjuder dig att ta ut lön nu, eftersom du fortsätter att styra av egen fri vilja.",
"##empire_service_tip##":"Sänd iväg trupper för att skydda",
"##dispatch_force##":"Sänd iväg undsättningsstyrka?",
"##dispatch_goods?##":"Sända iväg varor?",
"##legions##":"Legioner",
"##blessing_of_ceres_description##":"Förtjust över den uppmärksamhet som din stad visar henne förbättrar Ceres fruktbarheten hos din växande gröda.",
"##very_high_fire_risk##":"Mycket stor brandrisk",
"##collapse_available_damage_risk##":"Mycket stor risk för kollaps",
"##god_veryangry##":"Vredgade",
"##sldr_very_frightened##":"Mycket rädd",
"##god_quitepoor##":"Mycket dålig",
"##very_low_fire_risk##":"Mycket liten brandrisk",
"##some_defects_damage_risk##":"Mycket liten risk för kollaps",
"##sldr_very_bold##":"Mycket modig",
"##god_verypoor##":"Mycket dålig",
"##edu_poor##":"Mycket dålig",
"##non_cvrg##":"Mycket dålig",
"##god_charmed##":"Charmerade",
"##god_verygood##":"Mycket bra",
"##edu_awesome##":"Mycket bra",
"##statue_big_info##":"Monument över framstående medborgare och historiska händelser ger ett område bättre status. Folket är stolta över att ha statyer i grannskapet... och ju större desto bättre.",
"##barber_shop##":"Barberarsalong",
"##ovrm_barber##":"Barberare",
"##barbers##":"Barberarsalonger",
"##barber##":"Barberare",
"##wt_patrician##":"Patricier",
"##game_is_paused##":"Spelet pausat (Tryck P för att fortsätta)",
"##patients#":"patienter",
"##localization##":"LOKALISERING:",
"##send_to_city##":"Ge till staden",
"##give_money##":"Ge pengar",
"##send_money_to_city##":"Ge pengar till staden",
"##send_money##":"Donera dessa pengar till staden från dina personliga besparingar",
"##need_restart_for_apply_changes##":"Starta om spelet för att aktivera de nya inställningarna
",
"##goto##":"Gå till",
"##goto_empire_map##":"Gå till kartan över imperiet",
"##extm_troubles_tlp##":"Gå till problemområde.",
"##extm_reorient_map_to_north_tlp##":"Ändra visningen norrut",
"##egift_persian_carpets##":"Persiska mattor",
"##wn_picts##":"Pikter",
"##furniture_workshop_info##":"Snickarna vid snickeriet skapar fina möbler av virke. Medborgarna kan möblera sina villor och du kan handla med överskottet.",
"##empbutton_low_work##":"Fungerar dåligt. Tilldela fler människor till vår sektor",
"##poor_housing_discourages_migration##":"Dåliga bostäder motverkar invandring trots välståndet i staden",
"##sailing_to_city_docks##":"Seglar mot stadens lastkajer",
"##desirability_pretty_area##":"Detta land är ett eftertraktat område, vad gäller dina medborgare",
"##mission_win##":"Seger",
"##coast_caption##":"Kuster",
"##rotateRightBtnTooltip##":"Rotera panel medurs",
"##extm_rotate_map_clockwise_tlp##":"Rotera kartan medurs",
"##extm_rotate_map_counter_clockwise_tlp##":"Rotera kartan moturs",
"##rotateLeftBtnTooltip##":"Rotera panel moturs",
"##ovrm_damage##":"Skada
",
"##rioter_rampaging_accross_city##":"Kravaller i staden. De förstör och tar allt de kommer över.",
"##empire_tax##":"Tribut",
"##prepare_to_festival##":"Förbereder den kommande festivalen",
"##tooltip_full##":"Mushjälp - FULL",
"##tooltip_some##":"Mushjälp - DELVIS",
"##ovrm_fire##":"Brand",
"##fire##":"Brand",
"##donations##":"Donerat",
"##congratulations##":"Gratulerar",
"##tutorial_win_text##":"Gratulerar! Du har förstått grunderna på ett nöjsamt sätt. För att på bästa sätt fortsätta din utbildning, har jag ännu ett lindrigt uppdrag åt dig. Mot Brundisium!",
"##this_time_you_city_not_need_religion##":"Dina medborgare är ännu så länge upptagna med andra aspekter på stadslivet. I takt med att staden växer kommer de att vilja ha tillgång till ett stort Tempelutbud.",
"##freehouse_text##":"Ingen har så mycket som satt upp ett tält här ännu, fast immigranter kommer säkert att anlända inom kort om staden har tillgång till livsmedel och arbeten.",
"##cant_demolish_bridge_with_people##":"Kan inte förstöra bro med människor på",
"##have_no_requests##":"För närvarande har du inga meddelanden att läsa. I takt med att din stad växer, eller om kejsaren begär varor av dig, kommer meddelanden att visas här",
"##extm_show_bigpanel_tlp##":"Visa hela sidopanelen",
"##infobox_tooltip_help##":"Visa hjälpen för detta fönster",
"##show_prices##":"Visa priser",
"##btn_showprice_tooltip##":"Visar import-/exportpriser för alla varor, som anbefallt av Rom",
"##show##":"Evenemang",
"##leave_empire?##":"Lämna det Romerska Riket?",
"##coverage##":"Täckning i staden",
"##emw_buy##":"Inköp",
"##native_field##":"Ängmark
",
"##library_no_workers##":"Hyllorna i detta bibliotek är tomma, och värdelösa för lokalsamhället.",
"##granary_info##":"Fulla sädesmagasin är livsviktiga för att hålla folkets magar fyllda och för att attrahera nya medborgare. Ett sädesmagasin kan lagra säd, kött, grönsaker och frukt.",
"##fullscreen_on##":"Fullskärm",
"##deliver##":"Hämta varor",
"##no_dock_for_sea_trade_routes##":"GLÖM INTE! Denna nya handelsrutt över havet kräver byggnation av en handelshamn innan några fartyg kan anlända.",
"##gmenu_help##":"Hjälp",
"##help##":"Hjälp",
"##gmenu_shortkeys##":"Globala kortkommandon",
"##forum_information##":"En populär samlingsplats och eftertraktat samhällselement. Forum anställer även skatteindrivare och är livsviktiga för stadens skattkammare.",
"##dock_info##":"Hamnarbetarna hämtar varor som vi köper från lagerlokalen.",
"##dedicate_fectival_venus##":"Tillägna Venus en festival",
"##dedicate_fectival_mars##":"Tillägna Mars en festival",
"##dedicate_fectival_mercury##":"Tillägna Merkurius en festival",
"##dedicate_fectival_neptune##":"Tillägna Neptunus en festival",
"##dedicate_fectival_ceres##":"Tillägna Ceres en festival",
"##visit_military_advisor##":"Besök din militärrådgivare",
"##visit_chief_advisor##":"Besök din huvudrådgivare",
"##visit_imperial_advisor##":"Besök din imperierådgivare",
"##visit_health_advisor##":"Besök din hälsorådgivare",
"##visit_population_advisor##":"Besök din befolkningsrådgivare",
"##visit_education_advisor##":"Besök din utbildningsrådgivare",
"##visit_entertainment_advisor##":"Besök din underhållningsrådgivare",
"##visit_rating_advisor##":"Besök din ställningsrådgivare",
"##visit_religion_advisor##":"Besök din religionsrådgivare",
"##visit_trade_advisor##":"Besök din handelsrådgivare",
"##visit_labor_advisor##":"Besök din arbetsrådgivare",
"##visit_financial_advisor##":"Besök din finansrådgivare",
"##message_from_centurion##":"Från legion's centurion...",
"##dispatch_gift##":"Sänd en gåva",
"##dispatch_gift_title##":"Sänd gåva till kejsaren",
"##send_lavish_gift##":"Sänd en frikostig gåva",
"##send_modest_gift##":"Sänd en blygsam gåva",
"##send_generous_gift##":"Sänd en generös gåva",
"##engineer_low_entertainment##":"Efter en hård dags arbete vill jag se en bra pjäs eller strid. Det finns inte mycket chans till det i den här staden.",
"##barber_need_colloseum##":"Efter en dag med rakning och klippning vill jag se en trevlig lejonstrid. Men det går inte att uppbringa här.",
"##show_spots_of_city_troubles_tip##":"Växla mellan aktuella problemområden i staden",
"##barber_good_life##":"Rakning eller klippning, medborgare? Livet här är lätt att leva, inte sant?",
"##extm_road_tlp##":"Bygg vägar",
"##extm_housing_tlp##":"Bygg bostäder",
"##need_vines_farm##":"Bygg en vingård",
"##need_iron_mine##":"Bygg en järngruva",
"##need_timber_mill##":"Bygg en brädgård",
"##need_lionnursery##":"Bygg ett lejonhus för att arrangera djurtävlingar",
"##need_olive_farm##":"Bygg en olivodling",
"##need_actor_colony##":"Bygg en skådespelarkoloni för att sända skådespelare hit",
"##need_charioter_school##":"Bygg en skola för körsvenner för att se kapplöpningar",
"##colloseum_haveno_gladiatorpit##":"Bygg en gladiatorskola för att arrangera matcher här",
"##pottery##":"Krukor",
"##pottery_factory_stock##":"Krukor",
"##advchief_food_consumption##":"Matförbrukning",
"##sldr_shaken##":"Uppskakad",
"##cartPusher_normal_life##":"Allt verkar fungera bra här.",
"##engineer_average_life##":"Allt tycks fungera väl här.",
"##unhandled_key_8##":"Den här hopen tycks inte vara så lättskrämd.",
"##scholar_average_life##":"Den här staden verkar bra.",
"##taxCollector_average_life##":"Staden tycks fungera väl.",
"##favor_rating##":"Popularitetsställning",
"##valentia_preview_mission##":"Ståthållaren ställs inför olika hot och faror, och Iberierna utgör inte det minsta av dessa! De har inte för avsikt att ge upp Hispanien.",
"##win_syracusae_text##":"Bäste ståthållare, det var en lysande uppvisning. Du övertygade grekerna att överge sina planer för Syracusae vilket lägger hela Medelhavet för Roms fötter. Efter en sådan imponerande bragd kommer du aktivt att delta i framtida planer.",
"##rioter_say_1##":"Ståthållaren bryr sig uppenbarligen inte om mig, så jag tänker visa vad jag tycker om hans stad.",
"##festivals##":"Festivaler",
"##barracks_have_weapons_bad_workers##":"Med minimipersonal utbildar vi nya soldater mycket långsamt trots att vi har de vapen som krävs för att utbilda alla typer av soldater.",
"##city_warnings_on##":"Varningar: På",
"##city_warnings_off##":"Varningar: Av",
"##stop_granary_devastation##":"Sluta tömma sädesmagasin",
"##stop_warehouse_devastation##":"SLUTA tömma magasin",
"##desirability##":"Önskvärdhet",
"##ovrm_desirability##":"Prestige",
"##ovrm_crime##":"Brott",
"##wt_criminal##":"Brottsling",
"##prefect_low_entertainment##":"Brottslingarna jag tar får bättre underhållning än den här staden!",
"##advchief_crime##":"Brott",
"##layer_crime##":"Brott",
"##advchief_high_crime##":"Stor kriminalitet råder i staden",
"##advchief_which_crime##":"Brottsligheten håller på att bli ett problem.",
"##praetor##":"Praetor",
"##wt_prefect##":"Prefekt",
"##prefecture##":"Prefektur",
"##adve_prefectures##":"Prefekturer",
"##prefecture_info##":"Prefekturerna sänder prefekter till staden för att hålla fred, och för att bekämpa bränder. Ordning kan endast upprätthållas om prefekterna patrullerar staden.",
"##burning_ruins_info##":"Prefekterna kunde inte nå hit i tid för att rädda byggnaden. När elden har brunnit ut kommer endast spillror att finnas kvar på denna plats.",
"##engineer_high_workless##":"Jag har tur som har ett arbete i denna tid av arbetslöshet.",
"##romeGuard_high_workless##":"I dessa tider av arbetslöshet tackar jag gudarna att jag har jobb.",
"##city_under_rome_attack##":"De legioner från imperiet som närmar sig skrämmer dina invånare och förbättrar inte din fredsställning.",
"##city_zoom_on##":"Zoom: På",
"##city_zoom_off##":"Zoom: Av",
"##centurion_new_order_to_save_player##":"Nya order har just anlänt. Verkar som att Kjesaren har ändrat sig angående dig, och tacksamt ska jag återvända till Rom. Farväl...för denna gång.",
"##marketKid_say_3##":"Var hälsad! Jag bär korgen med mat till kvinnans marknad. Jag hoppas jag får bra med dricks!",
"##recruter_high_workless##":"Var hälsad! Har du sett hur hög arbetslösheten är?",
"##gladiator_gods_angry##":"Var hälsad, medborgare. Har du hört? Gudarna är vreda.",
"##gladiator_good_life##":"Var hälsad. Livet här är skönt att leva, inte sant?",
"##doctor_need_workers##":"Var hälsad! Det saknas många arbetare här.",
"##patrician_so_hungry##":"Hell! Vad tjänar rikedom till om det inte finns mat att köpa?",
"##wt_missioner_average_life##":"Var hälsad! Jag ser att det finns mycket att göra med att lära dessa barbarer fördelarna med Roms välvilja.",
"##missioner_high_barbarian_risk##":"Var hälsad! Min undervisning om Roms välvilja tycks tränga in hos dessa ganska skrämmande barbarer.",
"##engineer_good_life##":"Var hälsad! Är det inte en fantastisk stad?",
"##partician_good_life##":"Var hälsad. Staden sköts riktigt bra.",
"##taxCollector_good_life##":"Var hälsad! Detta är en mycket trevlig stad att bo i.",
"##priest_so_hungry##":"Var hälsad. Denna stad behöver omedelbart mer livsmedel.",
"##lionTamer_good_education##":"Var hälsad. Den här staden tycker vi om, inte sant, Leo?",
"##recruter_good_life##":"Var hälsad! Livet här är gott.",
"##recruter_normal_life##":"Var hälsad. Detta är en ganska bra stad.",
"##workers_yearly_wages_is##":"Beräknad årlig kostnad för",
"##accepting##":"Accepterar",
"##accept_goods##":"Acceptera varor",
"##may_collect_about##":"ger en avkastning på",
"##accept##":"Acceptera",
"##accept_promotion##":"Acceptera befordran",
"##accept_deity_status##":"Acceptera ställningen som kejsare!",
"##advemployer_panel_priority##":"prioritering",
"##fishing_wharf##":"Fiskehamn",
"##wharf##":"Fiskehamn",
"##docked_buying_selling_goods##":"Ligger vid kaj, köper och säljer varor",
"##migration_lack_tax##":"Höga skatter är ett problem",
"##migration_high_lack_workless##":"Hög arbetslöshet är ett problem",
"##low_wage_lack_migration##":"Låga löner är ett problem",
"##migration_low_food_stocks##":"Bristen på mat är ett problem",
"##ovrm_troubles##":"Problem",
"##new_festival##":"Anordna ny festival",
"##hold_venus_festival##":"Anordna festival för Venus",
"##hold_mars_festival##":"Anordna festival för Mars",
"##hold_mercury_festival##":"Anordna festival för Merkurius",
"##hold_neptune_festival##":"Anordna festival för Neptunus",
"##hold_ceres_festival##":"Anordna festival för Ceres",
"##arrange_festiable_for_this_god##":"Arrangera en festival till denna guds ära",
"##emw_sell##":"Försäljningar",
"##emw_sold##":"Sålt",
"##continue##":"Fortsätt",
"##mainmenu_continueplay##":"Fortsätt",
"##plname_continue##":"Fortsätt",
"##continue_2_years##":"Fortsätt att styra i 2 år till.",
"##continue_5_years##":"Fortsätt i 5 år till.",
"##operations_manager##":"Spelproducent",
"##industry_enabled##":"Industri är PÅ",
"##industry_disabled##":"Industri är AV",
"##adve_food##":"Livsmedelsproduktion",
"##rawm_production_complete_m##":"Produktionen är",
"##cursed_by_mars##":"Förbannad av Mars!",
"##proconsul##":"Proconsul",
"##procurator##":"Procurator",
"##line_formation_text##":"En enkel formation, som ger fördelar åt försvarstrupper.",
"##wt_rprotestor##":"Demonstrant",
"##senatepp_prsp_rating##":"Välstånd",
"##wndrt_prosperity##":"Välstånd",
"##percents##":"Ränta på",
"##month_from_last_festival##":"sedan senaste festivalen",
"##last_year##":"Förra året",
"##clear_land_caption##":"Tomt land",
"##engineer_gods_angry##":"Måtte gudarna vara mig nådiga. Det är inte mitt fel att ståthållaren hånar dem.",
"##wheat_farm##":"Veteodling",
"##warehouse_devastation_mode_text##":"Försöker sända gods till annan plats",
"##granary_devastation_mode_text##":"Försöker att sända mat till annan plats",
"##work##":"I bruk",
"##advemployer_panel_haveworkers##":"arbete",
"##abwrk_working##":"fungerar",
"##advemployer_panel_workers##":"arbetare",
"##unhandled_key_value_7##":"Fungerar med reducerad kapacitet. För få anställda har anlänt nyligen",
"##empbutton_simple_work##":"Fungerar, men fler arbetare skulle kunna tilldelas oss",
"##working_industry##":"fungerande industri i staden",
"##working_industries##":"fungerande industrier i staden",
"##forum_full_work##":"För närvarande arbetar våra indrivare med maximal effektivitet, och de är alltid ute och kontrollerar att alla förfallna skatter betalas in till staden.",
"##employee##":"Enhet",
"##employees##":"Enheter",
"##warehouseman##":"Magasinsman",
"##dock_bad_work##":"Vi har mycket få hamnarbetare så det kommer att ta lång tid att lasta och lossa de fartyg som anlöper hamnen.",
"##employers##":"Anställd arbetsstyrka",
"##healthadv_some_regions_need_hospital##":"Utvecklingen i vissa områden hålls tillbaka av för få sjukhus i staden. Nya sjukhus attraherar fler patricierklasser till staden.",
"##entertainment_short##":"Underhållning",
"##entertainmentBtnTooltip##":"Underhållning
",
"##adve_entertainment##":"Underhållning",
"##entertainment_advisor_title##":"Underhållning",
"##advchief_entertainment##":"Underhållning",
"##extm_entertainment_tlp##":"Underhållning",
"##entertainment##":"Underhållning",
"##ovrm_entertainments##":"Underhållning",
"##smallcurse_of_neptune_description##":"Neptunus är missnöjd med att du inte visar honom tillräcklig uppmärksamhet och frammanar en mindre storm.",
"##smallcurse_of_mars_description##":"Mars ogillar din brist på vördnad och sporrar ett antal missnöjda invånare att revoltera.",
"##god_wrathful##":"Rasande",
"##god_irriated##":"Sårade",
"##other##":"Diverse",
"##damage##":"Skador",
"##lawless_area##":"Ett laglöst område. Människorna är vettskrämda.",
"##loading_resources##":"Laddar tillgångar",
"##advemployer_panel_title##":"Arbetstilldelning",
"##smallcurse_of_ceres_description##":"Ceres är missnöjd med din brist på vördnad och ödelägger hela din skörd som en varning till dig.",
"##credit##":"Utgifter",
"##extm_clear_tlp##":"Röj marken",
"##reservoir##":"Reservoar",
"##need_connect_to_other_reservoir##":"Reservoir bör vara ansluten till vattnetskälla",
"##your_prosperity_raising##":"Din välståndsställning förbättras.",
"##wndrt_peace##":"Fredsställning",
"##peace_rating_text##":"Fredsställningen blir bättre för varje år utan upplopp eller invasioner som skadar egendom i städerna.",
"##rating##":"Ställning",
"##wnd_ratings_title##":"Ställning",
"##religion_advisor##":"Religiösa byggnader",
"##advchief_religion##":"Religion",
"##ovrm_religion##":"Religion",
"##religion##":"Religion",
"##religion_in_your_city_is_flourishing##":"Religionen i din stad blomstrar. Invånarnas olika religionsbehov uppfylls, och prästerna rapporterar att gudarna är nöjda.",
"##unhandled_key_value_6##":"Terrängen är bara ett av problemen du ställs inför här. Jämn mark är sällsynt, och det är svårt att transportera vatten till de högt belägna områdena.",
"##gmenu_file_restart##":"Starta om",
"##rome_gratitude_request_text##":"Rom tackar dig för din senaste sändning. Din lojalitet skall inte glömmas.",
"##your_favor_is_dropping_catch_it##":"Din popularitet i Rom minskar. Du måste fånga Caesars intresse på ett eller annat sätt!",
"##advemployer_panel_romepay##":"Rom betalar",
"##rome_raises_wages##":"Rom höjer lönerna",
"##try_reduce_your_high_salary##":"Rom tycker att din lön är för hög för din nuvarande ställning. Du borde sänka den lite.",
"##try_reduce_your_salary##":"Rom tycker att din lön är för hög för din nuvarande ställning. Det skulle vara bra om du sänkte den.",
"##rome_lowers_wages##":"Rom sänker lönerna",
"##roman_city##":"En romersk stad",
"##romechastener_attack_text##":"En romersk legion är inom sikte av staden. Detta är ett verkligen ett hot.",
"##rome_need_some_goods##":"Rom är i behov av följande varor. Var snäll och skicka dem så snabbt som möjligt.",
"##ovrm_risks##":"Risker",
"##beatifull_villa##":"Stor villa",
"##luxury_palace##":"Lyxpalats",
"##egift_lavish##":"Frikostig:",
"##lumber_mill_info##":"Såga virke för handel, eller till möbelverkstäderna. Patricierna vill ha möbler till sina villor, eller så kan du exportera det till dina handelspartners.",
"##collapsed_building_text##":"En byggnad har rasat. Dåligt underhåll av stadens ingenjörer av orsakat detta.",
"##fish##":"Fisk",
"##fishing_boat##":"Fiskebåt",
"##fishing_waters##":"Fiskevatten",
"##market##":"Marknad",
"##wt_marketLady##":"Marknadshandlare",
"##prosperity_lack_that_you_pay_less_rome##":"Att betala lägre löner än Rom ger din stad rykte att vara mindre blomstrande.",
"##marketBuyer_high_workless##":"Med denna höga arbetslöshet måste jag arbeta hårt för att behålla mitt jobb.",
"##factory_need_more_workers##":"Fungerar knappt. Tilldela fler människor till vår sektor",
"##partician_need_workers##":"Servicen blir lidande. Staden behöver fler arbetare.",
"##garden##":"Trädgårdar",
"##gardens_info##":"Trädgårdar förbättrar den lokala miljön.",
"##samnite_soldier##":"En samnitisk soldat",
"##wn_samnites##":"Samniter",
"##sarmizegetusa_title##":"Sarmizegetuza: en mycket farlig provins",
"##wt_taxCollector##":"Skatteindrivare",
"##lgn_pigs##":"Svinen",
"##free##":"ledig",
"##freehouse_caption##":"Ledig tomt",
"##north##":"Norr",
"##northBtnTooltip##":"Norr",
"##small_fest_description##":"En liten festival hölls denna kväll. Alla är tacksamma över detta avbrott i vardagen.",
"##theater_full_work##":"Denna teater sätter för närvarande upp pjäser med lokala aktörer, som vanligen drar stor publik.",
"##merchant_just_unloading_my_goods##":"Lagerlokalen lastar just av varor från mina djur.",
"##barracks_city_not_need_soldiers##":"Vi utbildar för närvarande inga rekryter eftersom vi inte har fått någon begäran från stadens fort eller torn om nya styrkor.",
"##dockers_taking_our_goods##":"Hamnarbetarna för våra varor till lagerlokalen nu.",
"##engineering_post_full_work##":"För närvarande har vi inga driftavbrott Våra ingenjörer är alltid ute och inspekterar och reparerar skador på stadens byggnader.",
"##well_haveno_houses_inarea##":"Denna brunn är överflödig för tillfället, eftersom det inte finns några hus inom dess serviceområde.",
"##merchant_little_busy_now##":"Jag är lite upptagen just nu.",
"##advemployer_panel_sector##":"Sektor",
"##seleucid_soldier##":"En selucidisk soldat",
"##wn_selecids##":"Selucider",
"##month_9_short##":"Sep",
"##senate_1##":"Senat",
"##extm_senate_tlp##":"Senat",
"##senate##":"Senat",
"##senate_1_info##":"Senatsbyggnaden är en av de attraktivaste byggnaderna i staden. Den ger anställning åt skatteindrivarna och inkomsterna från deras verksamhet förvaras här.",
"##warning_full##":"Varningar PÅ",
"##warning_some##":"Varningar AV",
"##sldh_health_strong##":"Stark",
"##sldr_badly_shaken##":"Mycket uppskakad",
"##rome_need_some_money##":"Jag ger dig härmed förmånen att tillhandahålla ytterligare medel för det goda i Rom. Skicka dem snart, och jag kommer att överväga att konstruera en staty i din ära.",
"##syracusae_title##":"Syracusae: en något farlig provins",
"##rock_caption##":"Klippor",
"##warehouse##":"Handelsmagasin",
"##stacking##":"Hamstrar",
"##stacking_resource##":"Hamstrar vara",
"##warehouses##":"Handelsmagasin",
"##city_have_goods_for_request##":"Dina lager rapporterar att du nu har tillräckligt av dessa varor för att uppfylla begäran från kejsaren.",
"##fountain_will_soon_be_hooked##":"Denna fontän väntar på att anslutas till det underjordiska rörledningsnätet.",
"##gmspdwnd_game_speed##":"Spelhastighet",
"##gmspdwnd_scroll_speed##":"Skrollningshastighet",
"##egift_modest##":"Blygsam:",
"##minimizeBtnTooltip##":"Göm panel",
"##hide_bigpanel##":"Göm sidopanelen, och utöka spelvyn",
"##sldh_health_sparse##":"Gles",
"##gladiator_low_entertainment##":"Tråkigt! Det säger alla om det här stället, trots mina tappra insatser. Staden behöver verkligen mer underhållning.",
"##too_close_to_enemy_troops##":"För nära fiendestyrkorna!",
"##unhandled_key_value_5##":"För få människor tilldelade av arbetsrådgivaren",
"##difficulty##":"Svårighetsgrad",
"##overlays##":"Översikt",
"##ovrm_text##":"Översikt",
"##sldr_daring##":"Djärv",
"##emperor_changed_title##":"Byte av kejsare",
"##bolt##":"Armborst",
"##taxСollector_low_tax_collected##":"Att driva in skatt från dessa hårt arbetande människor får mig nästan att gråta - men bara nästan!",
"##sldr_totally_distraught##":"Vettskrämd",
"##infobox_construction_comma_tip##":"TIPS: Använd komma och punkt för snabbflyttning genom dessa och andra objekt.",
"##trade_advisor##":"Handelsrådgivare",
"##advisors##":"Senat",
"##gmenu_advisors##":"Rådgivare",
"##soldier##":"Soldat",
"##soldiers_in_legion##":"Soldater i legion",
"##egift_soldier_from_pergamaum##":"En soldat från Pergamon",
"##soldiers##":"Soldater",
"##message##":"Meddelande",
"##no_warning_for_us##":"Vi har inga rapporter om hot",
"##advlegion_noalarm##":"Vi har inga rapporter om hot mot staden",
"##messages##":"Meddelanden",
"##extm_message_tlp##":"Meddelanden från dina skrivare",
"##scribe_messages_title##":"Meddelanden från dina skrivare",
"##nearby_building_negative_effect##":"En närliggande {0} har en försämrande effekt på efterfrågan till området. Försök att anlägga t ex trädgårdar, torg och statyer.",
"##advpopulation_text_census##":"Befolkningssammansättning efter ålder (år)",
"##advpopulation_text_society##":"Befolkningssammansättning efter inkomst",
"##savedlg_continue##":"Spara",
"##gmenu_file_save##":"Spara spel",
"##save_city##":"Spara spel",
"##save_map##":"Spara karta",
"##save_game_here##":"Spara det aktuella spelet till denna fil",
"##current_play_runs_for_another##":"Nuvarande pjäs spelas i ytterligare",
"##amphitheater_haveno_shows##":"Inga pjäser för närvarande",
"##special_orders##":"Specialorder",
"##demand##":"Krav",
"##middle_palace##":"Medelstort palats",
"##middle_insula##":"Medelstor Insulae",
"##middle_villa##":"Medelstor villa",
"##statue_middle##":"Medelstor staty",
"##tax_rate##":"Skattesatsen",
"##advlegion_window_title##":"Legionstatus",
"##become_trade_center##":"Utse till handelscentral",
"##wall##":"Mur",
"##wall_info##":"Murar skyddar värnlösa medborgare från barbarer. De kan bara motstå en viss grad av attacker, och tjockare murar klarar sig längre.",
"##fortification_info##":"Murar saktar ner fiendens framstöt mot en stad. Murar kan raseras. Tjockare murar är starkare och dessutom ges vaktposterna i anslutna torn möjlighet att patrullera dem.",
"##cost##":"Kostnad",
"##cost_2_open##":"Kostnad att öppna",
"##costs##":"kostnader",
"##wrath_of_venus_description##":"Tyvärr för dina olyckliga medborgare, Venus har inget annat val än att dela sin olycka, sprider sjukdom och elände hela folket.",
"##arrow##":"Pil",
"##ovrm_build##":"Byggnad",
"##buildings##":"Byggnation",
"##need_build_on_cleared_area##":"Måste byggas på avröjt land",
"##clay_pit_need_close_to_water##":"Bygg lertag nära vattnet",
"##timber_mill_need_trees##":"Bygg brädgård intill träden",
"##build_markets_to_distribute_food##":"Bygg marknader för att distribuera maten som lagrats här",
"##farm_need_farmland##":"Bygg jordbruk på jordbruksmark (leta efter gult gräs)",
"##students##":"i högskoleålder.",
"##egift_chest_of_sapphire##":"En kista med safirer",
"##god_happy##":"Glada",
"##bldm_raw_material##":"Råmaterial",
"##tarentum_title##":"Tarente: une petite province dangereuse",
"##tarentum_slightly_dangerous_province##":"Tarentum: en inte helt ofarlig provins",
"##tarraco_title##":"Tarraco: en fredlig provins",
"##tarsus_title##":"Tarsus: en mestadels fredlig provins",
"##theater##":"Teater",
"##ovrm_theater##":"Teatrar",
"##theaters##":"Teatrar",
"##theater_need_actors##":"Teatrarna och amfiteatrarna söker alltid efter nya talanger.",
"##population_tooltip##":"Befolkningsmängd",
"##finance_advisor##":"Stadens kapital",
"##scrw_subject##":"Ämne",
"##tingis_title##":"Tingis: en farlig provins",
"##your_province_quiet_and_secure##":"Din provins lugna och säkra tillvaro har blivit legendarisk. Andra ståthållare planerar förmodligen att dra sig tillbaka hit!",
"##mediolanum_win_text##":"Att Hannibal kunde korsa Alperna med sina elefanter var häpnadsväckande. Att Mediolanum skulle blomstra trots hans attacker är ett mirakel. Din framgång vände lyckan i det puniska kriget till Roms fördel. Hela Rom tackar dig.",
"##emperor_send_money_to_you_nearest_time##":"Det faktum att kejsaren nyligen måste ingripa för att rädda dig skadar allvarligt din stads rykte om välstånd.",
"##warehouse_info##":"Varor som produceras för handel kräver magasinering. Karavaner besöker handelsmagasinen för att köpa och sälja varor och handelshamnar får sitt gods från intilliggande magasin.",
"##cartPusher_low_entertainment##":"...vagnar. Det är mer underhållande än resten av den här staden.",
"##mercury_desc##":"Handel",
"##trade##":"Handel",
"##small_mercury_temple_info##":"Handelsmännen dyrkar Merkurius för att skydda sina varor. Om Merkurius vrede väcks sätts allas vinst på spel.",
"##dock_about##":"Handelsskepp från hela riket lägger till här för att leverera importvaror och hämta exportvaror. Du kan inte bedriva sjöhandel utan en handelshamn.",
"##no_working_dock##":"Varningar",
"##trading_city##":"Handelsstad",
"##trade_caravan_from##":"Köpmannakaravan från",
"##trade_ship_from##":"Handelsskepp från",
"##trade_center##":"Handelscentral",
"##trading_goods##":"Byter varor",
"##exit_point##":"Utträdespunkt",
"##grass##":"Gräs",
"##imperial_request##":"Kejserlig begäran",
"##requierd##":"Behov",
"##demands_3_religion##":"Krav på tillgång till en tredje religion",
"##need_population##":"krävs)",
"##crack##":"Spricka",
"##rift_info##":"Sprickor i marken",
"##triumphal_arch##":"Triumfbåge",
"##labor##":"Arbetskraft",
"##land_trade_problem_title##":"Problem med landhandeln",
"##egift_troupe_preforming_slaves##":"En grupp uppträdande slavar",
"##wt_indigene##":"Inföding",
"##wn_indigene##":"Infödingar",
"##recruter_so_hungry##":"Kan du avvara lite bröd? Jag har inte ätit på så länge.",
"##nomoney_for_gift_text##":"Du har inte tillräcklig med personliga besparingar för att kunna betala en gåva till kejsaren. Försök att betala dig själv högre lön!",
"##legionadv_no_legions##":"Du har inga legioner att leda. Du måste först bygga ett fort",
"##have_no_legions##":"Du har inga legioner att sända",
"##city_has_runout_debt##":"Din stad har inga pengar kvar. Caesar har gått med på att ge dig mer, men han kommer inte vara så generös nästa gång. Exportera varor för att generera mer inkomst till din stad.",
"##healthadv_noproblem_small_city##":"Din lilla bosättning har ännu inga hälsoproblem att rapportera.",
"##city_has_runout_money##":"Din stad har inga pengar kvar. Caesar har gått med på att ge dig mer, men han kommer inte vara så generös nästa gång. Exportera varor för att generera mer inkomst till din stad.",
"##emperor_favour_10##":"Kejsaren är fundersam vad gäller dig.",
"##tower_have_workers_no_soldiers##":"Vi har underhållspersonal, men vi behöver trupper från en förläggning för att försvara staden.",
"##engineering_post_need_some_workers##":"Det tar en eller två dagar innan våra utarbetade ingenjörer är tillbaka på gatorna.",
"##barracks_have_weapons_slow_workers##":"Vi är underbemannade och utbildar nya soldater långsamt, men vi har de vapen som krävs för att utbilda alla typer av soldater.",
"##lion_pit_patrly_workers##":"Vi har bara halva personalstyrkan, och kan därför endast leverera ett lejon under nästa månad.",
"##actorColony_patrly_workers##":"Vi har bara halva personalstyrkan, och kan därför endast utbilda en skådespelare under nästa månad.",
"##gladiator_pit_patrly_workers##":"Vi har bara halva personalstyrkan, och kan därför endast utbilda en gladiator under nästa månad.",
"##charioteer_school_patrly_workers##":"Vi har bara halva personalstyrkan, och kan därför endast tillverka en vagn under nästa månad.",
"##forum_patrly_workers##":"Vi är underbemannade och måste vänta en vecka innan våra indrivare är tillbaka i tjänst.",
"##dock_need_some_workers##":"Vi är underbemannade och därför kommer det att ta lite längre tid än vanligt att lasta och lossa de fartyg som anlöper hamnen.",
"##recruter_gods_angry7##":"Vi har problem! Gudarna är förargade på oss.",
"##prefecture_slow_work##":"Vi har alldeles för få prefekter. Det händer att inga prefekter lämnar stationen på upp till två veckor åt gången.",
"##forum_need_some_workers##":"Vi har korta avbrott i verksamheten, ungefär en dag eller två, innan våra indrivare är tillbaka på gatorna igen.",
"##unhandled_key_value_4##":"Med så få anställda tar det oss en månad mellan varje gång vi sänder ut indrivare.",
"##education_have_academy_access##":"Detta hus har tillgång till högskola",
"##awesome_amphitheater_access##":"Detta hus har tillgång till amfiteater",
"##baths_full_access##":"Detta hus har tillgång till badhus",
"##library_full_access##":"Detta hus har tillgång till bibliotek",
"##hospital_full_access##":"Detta hus har tillgång till sjukhus",
"##hippodrome_full_access##":"Detta hus har tillgång till hippodrom",
"##awesome_doctor_access##":"Detta hus har tillgång till en klinik",
"##awesome_colloseum_access##":"Detta hus har tillgång till colosseum",
"##religion_access_full##":"Detta hus har tillgång till ett orakel, och till tempel för alla gudar",
"##barber_full_access##":"Detta hus har tillgång till barberare",
"##theater_full_access##":"Detta hus har tillgång till teater",
"##religion_access_5_temple##":"Detta hus har tillgång till tempel för alla gudarna",
"##religion_access_2_temple##":"Detta hus har tillgång till tempel för 2 olika gudar",
"##religion_access_3_temple##":"Detta hus har tillgång till tempel för 3 olika gudar",
"##religion_access_4_temple##":"Detta hus har tillgång till tempel för 4 olika gudar",
"##religion_access_1_temple##":"Detta hus har endast tillgång till ett tempel för en enda gud",
"##school_full_access##":"Detta hus har tillgång till skola",
"##education_full_access##":"Detta hus har tillgång till skola, bibliotek och högskola",
"##education_have_school_or_library_access##":"Detta hus har tillgång till skola eller bibliotek",
"##education_have_school_library_access##":"Detta hus har tillgång till skola och bibliotek",
"##no_academy_access##":"Detta hus har inte tillgång till en högskola",
"##amphitheater_no_access##":"Detta hus har inte tillgång till en amfiteater",
"##library_no_access##":"Detta hus har inte tillgång till bibliotek",
"##hospital_no_access##":"Detta hus har inte tillgång till ett sjukhus",
"##hippodrome_no_access##":"Detta hus har inte tillgång till hippodromen",
"##doctor_no_access##":"Detta hus har inte tillgång till en klinik",
"##colosseum_no_access##":"Detta hus har ingen tillgång till ett colosseum",
"##barber_no_access##":"Detta hus har inte tillgång till en barberare",
"##bath_no_access##":"Detta hus har inte tillgång till ett fungerande badhus",
"##theater_no_access##":"Detta hus har inte tillgång till en teater",
"##religion_no_access##":"Detta hus har inte tillgång till några tempel eller orakel",
"##school_no_access##":"Detta hus har inte tillgång till någon skola",
"##education_have_no_access##":"Detta hus har ingen grundläggande tillgång till skolor eller bibliotek",
"##house_no_troubles_with_food##":"Detta hus har inget problem med att skaffa den mat som krävs för att överleva",
"##awesome_entertainment_access##":"Denna boning har tillgång till flera platser för underhållning",
"##9_entertainment_access##":"Denna boning har tillgång till all underhållning som kan önskas",
"##2_entertainment_access##":"Denna boning har viss tillgång till underhållning",
"##1_entertainment_access##":"Denna boning har knappt tillgång till underhållning",
"##0_entertainment_access##":"Denna boning har inte tillgång till underhållning överhuvudtaget",
"##5_entertainment_access##":"Denna boning har begränsad tillgång till underhållning",
"##8_entertainment_access##":"Denna boning har utmärkt tillgång till underhållning",
"##3_entertainment_access##":"Denna boning har mycket begränsad tillgång till underhållning",
"##7_entertainment_access##":"Denna boning har mycket god tillgång till underhållning",
"##4_entertainment_access##":"Denna boning har rimlig tillgång till underhållning",
"##6_entertainment_access##":"Denna boning har god tillgång till underhållning",
"##trouble_most_damage##":"Denna byggnad har många strukturella brister och sprickor",
"##very_low_damage_risk##":"Denna byggnad har vissa strukturella brister",
"##some_low_fire_risk##":"Denna byggnad utgör en försumbar brandrisk",
"##trouble_some_damage##":"Denna byggnad löper försumbar risk att kollapsa",
"##middle_file_risk##":"Denna byggnad har en viss brandrisk",
"##trouble_have_damage##":"Denna byggnad löper en liten risk att kollapsa",
"##fired##":"Avskedad!",
"##distant_city##":"En avlägsen stad",
"##delete##":"Radera",
"##delete_game##":"Radera spelet",
"##delete_object##":"Radera objekt",
"##delete_this_message##":"Radera detta meddelande",
"##granary_orders##":"Instruktioner sädesmagasin",
"##warehouse_orders##":"Instruktioner handelsmagasin",
"##access_ramp##":"Åtkomstramp",
"##wt_lion_tamer##":"Lejontämjare",
"##destroy_bridge##":"Förstör en bro
",
"##destroy_fort##":"Förstör ett fort",
"##poor_city_mood_lack_migration##":"Stämningen i staden förhindrar immigration",
"##adve_administration_religion##":"Styrelse/Religion",
"##doctor_high_workless##":"Arbetslösheten är mycket hög. Jag funderar på att ge mig av.",
"##cartPusher_high_workless##":"...min fru har slutat tjata om att jag ska skaffa mig ett nytt arbete.",
"##citizen_high_workless10##":"Arbetslösheten är så hög att hela staden mår dåligt.",
"##advchief_health_simple_clinic##":"Stadens hälsosituation är mindre bra",
"##advchief_health_simple##":"Stadens hälsosituation är inte bra, se till att dina medborgare har mat och kliniker.",
"##advchief_health_bad##":"Stadens hälsosituation är dålig",
"##advchief_health_bad_clinic##":"Stadens hälsosituation är dålig, dina överansträngda läkare fruktar en dödlig epidemi.",
"##priority_level##":"Prioritetsnivå",
"##adve_water##":"Vattenförsörjning",
"##wage_level_tip##":"Fastställ en lönenivå (ditt folk kommer att jämföra denna med lönerna i Rom)",
"##set_amount_to_donate##":"Fastställ summa att donera",
"##wt_teacher##":"Lärare",
"##unhandled_key_value_3##":"Sårbar romersk stad",
"##file##":"Arkiv",
"##month_2_short##":"Feb",
"##wt_surgeon##":"Kirurg",
"##farm##":"Lantbruk",
"##bldm_farm##":"Jordbruk",
"##advchief_finance##":"Finanser",
"##finance_title##":"Finanser",
"##finances##":"Finanser",
"##fountain##":"Fontän",
"##fort##":"Fort",
"##fort_legionaries##":"Legionärfort",
"##fort_info##":"Ett romerskt fort rekryterar soldater från förläggningar. Lägga till en militärhögskola skulle ge trupper med bättre utbildning.",
"##forum##":"Forum",
"##fig_farm##":"Fruktodling",
"##fruit##":"Frukt",
"##fig_farm_info##":"Frukt är en viktig del av den balanserad diet som ditt folk behöver för hälsa och glädje. I sädesmagasinen lagras frukt för lokal konsumtion, och i handelsmagasinen förvaras överskottet för export.",
"##native_hut##":"Infödingshydda",
"##god_good##":"Bra",
"##hospital_info##":"Även om ingen vill bo i närheten av dem, räddar sjukhus liv. Staden borde ha tillräckligt med sängplatser för alla sina invånare.",
"##small_venus_temple##":"Venustempel",
"##small_mars_temple##":"Marstempel",
"##small_mercury_temple##":"Merkuriustempel",
"##small_neptune_temple##":"Neptunustempel",
"##small_ceres_temple##":"Cerestempel",
"##temples##":"Tempel",
"##extm_temples_tlp##":"Tempel",
"##units_in_stock##":"Lagrar",
"##qty_stacked_in_city_warehouse##":"förvaras i stadens handelsmagasin",
"##сaesar##":"Caesar",
"##caesar_assign_new_title##":"Caesar har befordrat dig till graden",
"##emperoradv_caesar_has_high_respect_for_you##":"Caesar respekterar dig mer än någon annan ståthållare någonsin!",
"##mission_wnd_targets_title##":"Mål",
"##buy_price##":"Köparna betalar",
"##sell_price##":"Säljarna får",
"##native_center##":"Inhemskt centrum",
"##rome_prices##":"Priser fastställs av Rom",
"##god_ceres_short##":"Ceres",
"##ceres_goodmood_info##":"Ceres skänker fruktsamhet åt jorden, och får plantorna att växa. Blidka henne, eller bered dig på hungersnöd.",
"##smallcurse_of_ceres_title##":"Ceres är upprörd",
"##baths_info##":"Civiliserade människor badar minst en gång om dagen. Utöver bättre hälsa utgör baden även en önskvärd träffpunkt med olika rekreativa aktiviteter.",
"##wt_endeavor##":"Endeavor",
"##wt_romeGuard##":"Vaktpost",
"##money_stolen_text##":"Fortfarande frustrerad, några invånare har börjat stjäla. De mer laglydiga invånarena har börjat prata om att flytta. Handla nu för att förbättra humöret på dem.",
"####unhandled_key_value_2##":"Vissa av våra trupper behövs på annan plats i riket",
"##person##":"denarer",
"##more_people##":"Anställda",
"##more_person##":"Anställd",
"##trees_and_forest_text##":"Träden kan inte forceras, men de kan röjas undan. De är livsviktiga för skogsindustrin, brädgårdar måste ligga nära träden för att producera timmer.",
"##rock_text##":"Klipporna kan inte forceras eller röjas undan. Marmor- och malmbrott fungerar bara om de uppförs nära klippor.",
"##profit##":"Nettoflöde in/ut",
"##defensive_formation_text##":"En mycket defensiv formation. Nästan omöjlig att penetreras av missiler.",
"##overall_city_become_a_sleepy_province##":"Detta är på det hela taget en provins med få verkliga hot - precis så som invånarna vill ha det!",
"##cartPusher_so_hungry##":"...dagen kräver styrka. Hur ska en vagndragare kunna arbeta utan mat?",
"##school##":"Skola",
"##actorColony##":"Skådespelarkoloni",
"##chatioteer_school##":"Skola för körsvenner",
"##chatiotSchool##":"Skola för körsvenner",
"##gladiator_pit##":"Gladiatorskola",
"##gladiatorSchool##":"Gladiatorskola",
"##ovrm_school##":"Skola",
"##schools##":"Skolor",
"##scholar##":"Skolbarn",
"##scholars##":"i skolålder",
"##roadBlock##":"Vägstopp",
"##warehouse_no_workers##":"Endast minimibemanning. Kommer ej att sända eller ta emot varor",
"##egift_generous##":"Generös:",
"##minimap_tooltip##":"Klicka på denna översiktskarta för att flytta till avlägsna delar av din stad",
"##click_item_for_start_trade##":"Klicka på en vara",
"##click_on_city_for_info##":"Klicka på en stad för att få information",
"##click_on_rating_for_info##":"Klicka på en stad för att få information",
"##right_click_to_exit##":"Högerklicka för att avsluta",
"##left_click_open_right_erase##":"Vänsterklicka på ett meddelande för att läsa. Högerklicka för att radera.",
"##aedile##":"Edil",
"##extm_comerce_tlp##":"Handel",
"##commerce##":"Handel",
"##export##":"Export",
"##tarraco_win_text##":"Tarracos livsmedelsexport hjälpte imperiet att överleva en svår period. Medborgarna är skyldiga dig för sina liv och ståthållarna sina arbeten. Skördarna blir nu normala igen och jag vill använda dina talanger inom ett nytt område.",
"##exports_over##":"Exportera vara över",
"##trade_btn_export_text##":"Exportera vara över",
"##wt_emigrant##":"Emigrant",
"##emigrant##":"Emigrant",
"##academy_no_workers##":"Denna högskola används inte, och är därför värdelös för lokalsamhället.",
"##academy_full_work##":"Denna högskola används, och ungdomarna i stadsdelen lär sig sociala färdigheter.",
"##library_full_work##":"Detta bibliotek används. Dess hyllor är fyllda med skriftrullar med lärdom.",
"##hospital_no_workers##":"Detta sjukhus används inte, och är därför värdelöst för lokalsamhället.",
"##hospital_full_work##":"Detta sjukhus används, och betjänar lokalsamhället.",
"##wine_workshops_patrly_workers##":"Denna vingård utnyttjar inte full kapacitet. Vinproduktionen något långsammare än vad den borde vara.",
"##road_from_rome##":"Detta är vägen till Rom. Immigranterna anländer från denna punkt. Därför är det viktigt att vägen hålls öppen. Även köpmän passerar genom din provins längs denna kejserliga huvudväg.",
"##this_lawab_province_become_very_peacefull##":"Detta är en laglydig provins som med tiden kan bli mycket fredlig.",
"##clinic_no_workers##":"Denna klinik används inte, och är därför värdelös för lokalsamhället.",
"##clinic_full_work##":"Denna klinik används, och betjänar lokalsamhället.",
"##marketKid_say_2##":"Korgen tar kål på mig. Jag bryr mig inte om vem som behöver maten, det borde finnas en lag mot barnarbete.",
"##lumber_mill_need_some_workers##":"Denna brädgård arbetar inte med maximal kapacitet. Som resultat kommer timmerproduktionen att bli något långsammare.",
"##wine_workshop_need_resource##":"Denna vingård kan inte producera vin förrän den får en leverans av druvor från ett magasin eller en druvodling.",
"##oil_workshop_need_resource##":"Denna olivpress kommer inte att producera olja utan leverans av oliver, från ett magasin eller från en lantgård.",
"##weapons_workshop_patrly_workers##":"Denna smedja utnyttjas inte till maximal kapacitet. Vapenproduktionen kommer att gå något långsammare än vad den borde.",
"##pottery_workshop_patrly_workers##":"Detta krukmakeri utnyttjar inte maximal kapacitet. Som resultat kommer krukproduktionen att gå långsammare.",
"##barber_no_workers##":"Denna barberarlokal används inte, och är därför värdelös för lokalsamhället.",
"##barber_full_work##":"Denna barberarlokal används, och ortsbefolkningen är vältrimmad.",
"##nativeCenter_info##":"Mötesplatsen för den lokalbefolkning som kommer hit för att byteshandla med enkla handelsvaror. Om styresmannen bara kunde lära sig några ord på latin...",
"##province_has_peace_a_short_time##":"Denna provins har haft fred en kort tid, men dina invånare känner sig fortfarande inte helt säkra. Fler fredsår kommer att förbättra detta.",
"##trouble_farm_was_blighted_by_locust##":"Jordbrukets marker har skadats av gräshoppssvärmarna, återhämtningen kommer att ta tid.",
"##vegetable_farm_patrly_workers##":"Denna lantgård utnyttjar inte maximal kapacitet. Därför kommer grönsaksproduktionen att gå något långsammare.",
"##fig_farm_patrly_workers##":"Denna fruktträdgård utnyttjar inte maximal kapacitet. Som resultat kommer fruktproduktionen att gå långsammare.",
"##meat_farm_patrly_workers##":"Denna farm arbetar inte med maximal kapacitet. Som resultat kommer köttproduktionen att bli något mindre.",
"##olive_farm_need_some_workers##":"Denna lund utnyttjar inte maximal kapacitet. Olivproduktionen kan bli bättre med fler arbetare.",
"##wheat_farm_patrly_workers##":"Denna lantgård arbetar under sin maximala kapacitet. Fler arbetare skulle öka produktiviteten.",
"##school_no_workers##":"Denna skola används inte, och är värdelös för lokalsamhället.",
"##actorColony_no_workers##":"Denna koloni är övergiven. Utan tillgång till mentorer kan inga nya skådespelare utbildas.",
"##school_full_work##":"Denna skola används, och barnen i stadsdelen är läskunniga och vältaliga.",
"##population_milestone##":"Populations milstolpe",
"##baths_no_workers##":"Detta badhus används inte, och är därför värdelöst för lokalsamhället.",
"##baths_full_work##":"Detta badhus används, besökarna blir rena och avslappnade.",
"##baths_need_reservoir##":"Detta badhus behöver en rörledning till en reservoar.",
"##taxCollector_very_little_tax##":"Dessa hus betalar så lite skatt att det är slöseri med tiden.",
"##marketBuyer_return##":"Dessa korgar är så tunga! Jag har med mig färska varor till min marknad.",
"##nativeField_info##":"Vissa primitiva grödor, som förser lokalbefolkningen med en grundläggande källa till livsmedel.",
"##engineer_have_trouble_buildings##":"Dessa byggnader är i dåligt skick. Jag kom precis i rätt tid.",
"##collapsed_ruins_info##":"Dessa spillror av gamla byggnader gör marken mindre åtråvärd.",
"##these_rift_info##":"Dessa klyftor har orsakats av jordbävningar. De kan inte passeras eller fyllas.",
"##these_goods_import_only##":"Dessa varor finns endast tillgängliga via import",
"##marketBuyer_gods_angry##":"Detta är en hednisk plats. Ståthållaren har ingen respekt för gudarna.",
"##citizen_gods_angry##":"Detta är en hednisk stad. Den behöver fler tempel.",
"##cartSupplier_good_life##":"Detta är en magnifik stad.",
"##triumphal_arch_info##":"Detta magnifika byggnadsverk är tillägnat Roms historiska segrar över sina fiender. Inget kan ge högre status.",
"##inland_lake_text##":"Denna insjö saknar kontakt med havet",
"##priest_average_life##":"Denna stad är en hygglig plats att bo på.",
"##road_to_distant_region##":"Detta är den väg som leder till rikets utposter. Det är en kejserlig huvudväg, som måste hållas öppen längs hela sin sträckning.",
"##very_low_crime_risk##":"Detta är en mycket laglydig stadsdel, ingen brottslighet alls",
"##doctor_average_life##":"Detta är en fantastisk stad.",
"##trouble_most_fire##":"Denna byggnad är en brandfara",
"##trouble_low_fire_risk##":"Denna byggnad har ingen brandrisk",
"##no_space_for_evolve##":"Denna boning skulle kunna få ännu högre status om den hade mer utrymme att expandera.",
"##moment_fire_risk##":"Denna byggnad kan fatta eld när som helst!",
"##trouble_some_fire##":"Denna byggnad har brandrisk",
"##trouble_no_damage##":"Denna byggnad är i perfekt strukturellt skick",
"##very_high_damage_risk##":"Denna byggnad är ostadig, och kommer sannolikt att falla samman snart",
"##trouble_need_road_access##":"Denna byggnad kräver åtkomst till väg",
"##house_evolves_at##":"Denna boning kommer snart att utvecklas och få bättre status, som ett resultat av de förbättrade lokala villkoren.",
"##trouble_too_far_from_water##":"Denna byggnad är inte intill vatten!",
"##peaceful_crime_risk##":"Detta är en fridfull stadsdel.",
"##prefect_good_life##":"Detta är en underbar plats att bo på.",
"##this_province_feels_peaceful##":"Denna provins känns förhållandevis säker, en känsla som kan förbättras med tiden.",
"##garden_info##":"Denna trevliga plats skänker medborgarna avkoppling från stadens buller, värme och smuts genom en sval oas av grönska. Alla vill ha en trädgård intill sitt hus.",
"##this_is_ruins##":"Detta är spillrorna från byggnaden som nämns ovan. Förfallna platser gör inte att området ser vackrare ut.",
"##averange_crime_risk##":"Detta är ett område med hög brottslighet. De boende är missnöjda, och gatorna är farliga",
"##few_crime_risk##":"Detta är ett område med låg brottslighet, men vissa boende har klagat",
"##lionTamer_good_life##":"Nu har du din chans, Leo. Duktigt lejon.",
"##gladiator_need_workers##":"Det är hemskt. Jag har aldrig sett så många lediga jobb.",
"##cartSupplier_average_life##":"Det här är en bra stad. Folk tycker om att bo här.",
"##oil_workshop_patrly_workers##":"Denna olivpress är underbemannad och producerar oljan mycket långsammare än vad den borde.",
"##taxCollector_need_workers##":"Den här staden behöver fler arbetare och det genast.",
"##citizen_need_workers3##":"Staden lider stor brist på arbetare.",
"##citizen_need_workers5##":"Staden behöver fler arbetare!",
"##priest_need_workers##":"Detta ställe behöver många fler arbetare.",
"##romeGuard_need_workers##":"Den här staden behöver många fler arbetare.",
"##lionTamer_need_workers##":"Den här staden behöver mer arbetskraft. Jag undrar om jag kan träna Leo att arbeta mer?",
"##need_grape##":"Denna byggnad kräver druvor",
"##building_need_road_access##":"Denna byggnad behöver tillgång till väg",
"##need_clay_pit##":"Denna byggnad kräver lera",
"##trouble_need_timber##":"Denna byggnad kräver timmer",
"##need_iron_for_work##":"Denna byggnad kräver järnmalm",
"##trouble_need_olive##":"Denna byggnad kräver oliver",
"##aqueduct_no_water##":"Denna akvedukt transporterar inte vatten mellan reservoarer eftersom den saknar vattenkälla.",
"##aqueduct_work##":"Denna akvedukt transporterar vatten mellan reservoarer.",
"##amphitheater_have_never_show##":"Denna amfiteater har sällan några föreställningar. Den behöver skådespelare och gladiatorer.",
"##amphitheater_full_work##":"Denna amfiteater erbjuder sitt samhälle både intressant gladiatorkamp och pjäser med lokala skådespelare.",
"##amphitheater_have_only_battles##":"Denna amfiteater erbjuder gladiatorkamp som förströelse. Den söker skådespelare för att sätta upp några pjäser.",
"##amphitheater_no_workers##":"Denna amfiteater är stängd. Den har inga anställda, och erbjuder ingen förströelse åt det lokala samhället.",
"##amphitheater_have_only_shows##":"Denna amfiteater sätter upp pjäser med lokala aktörer. Den kan attrahera större publik om den även har gladiatorer.",
"##vinard_patrly_workers##":"Denna odling utnyttjar inte maximal kapacitet. Som resultat kommer druvproduktionen att bli mindre.",
"##engineer_need_workers##":"Staden skulle fungera bättre om det fanns nog med arbetare.",
"##citizen_good_education##":"Den här staden är mer kultiverad än någon annan i riket!",
"##prefect_need_workers##":"Denna stad är i desperat behov av arbetare!",
"##teacher_good_life##":"Staden får full pott. Det är en underbar plats.",
"##scholar_good_life##":"Den här staden är fantastisk.",
"##actor_good_life##":"Den här staden är inte så illa.",
"##doctor_low_entertainment##":"Staden är så trist att mina patienter frågar om jag kan bota kronisk uttråkning!",
"##teacher_low_entertainment##":"Staden är så tråkig! Den behöver mer underhållning.",
"##scholar_low_entertainment##":"Staden är så tråkig. Jag vill se fler föreställningar.",
"##priest_low_entertainment##":"Denna stad är så tråkig. Även en präst tycker om gladiatorspel då och då.",
"##marketBuyer_average_life##":"Denna stad är egentligen inte så illa.",
"##cartPusher_good_life##":"Stad som stad... Den här verkar rätt bra.",
"##house_not_registered_for_taxes##":"Detta hus befinner sig i en region utan skatteadministration, och betalar därför ingen skatt",
"##missing_entertainment##":"Detta hus kan inte utvecklas, eftersom det inte finns någon underhållning i området.",
"##missing_entertainment_amph##":"Detta hus kan inte utvecklas, eftersom det knappt finns någon underhållning i området.",
"##missing_entertainment_also##":"Detta hus kan inte utvecklas, eftersom det inte finns tillräckligt med underhållning i området.",
"##missing_library##":"Detta hus kan inte utvecklas, eftersom dess tillgång till utbildning måste förbättras genom tillgång till ett bibliotek.",
"##missing_school##":"Detta hus kan inte utvecklas, eftersom dess tillgång till utbildning måste förbättras genom tillgång till en skola.",
"##missing_college##":"Detta hus kan inte utvecklas, eftersom dess redan utmärkta tillgång till utbildning måste förbättras genom tillgång till en högskola.",
"##missing_second_food##":"Detta hus kan inte utvecklas, eftersom det krävs en till typ av livsmedel, som levereras från en lokal marknad, för att förmå mer välbärgade att flytta in.",
"##missing_third_food##":"Detta hus kan inte utvecklas, eftersom det krävs en tredje typ av livsmedel, som levereras från en lokal marknad, för att förmå patricierklasserna att flytta in.",
"##missing_hospital##":"Detta hus kan inte utvecklas, eftersom det vill ha bättre möjligheter till sjukvård. Klinikernas täckning är bra men det saknas lokal tillgång till ett sjukhus.",
"##missing_doctor##":"Detta hus kan inte utvecklas, eftersom det vill ha bättre möjligheter till sjukvård. Det finns lokal tillgång till ett sjukhus men det behövs en klinik i närheten.",
"##missing_food##":"Detta hus kan inte utvecklas, eftersom det måste ha leveranser av livsmedel från en lokal marknad.",
"##missing_entertainment_patrician##":"Detta hus kan inte utvecklas, eftersom det visserligen finns utmärkt underhållning i området, men det är trångt och utbudet är inte tillräckligt varierat för de kräsna patricierna.",
"##missing_entertainment_colloseum##":"Detta hus kan inte utvecklas, eftersom det visserligen finns viss underhållning i området, men inte tillräckligt.",
"##missing_third_religion##":"Detta hus kan inte utvecklas, eftersom det endast har tillgång till tempel för två gudar. I takt med att dess invånare kommer upp sig i världen kommer de att vilja ägna mer tid åt att tillbe andra gudar.",
"##missing_second_religion##":"Detta hus kan inte utvecklas, eftersom det endast har tillgång till tempel för en enda gud. I takt med att dess invånare kommer upp sig i världen kommer de att vilja ägna mer tid åt att tillbe andra gudar.",
"##missing_water##":"Detta hus kan inte utvecklas, eftersom det inte har tillgång till ens den mest primitiva vattenförsörjning.",
"##missing_market##":"Detta hus kan inte utvecklas, eftersom det inte har tillgång till en lokal marknad.",
"##missing_bath##":"Detta hus kan inte utvecklas, eftersom det inte har tillgång till ett lokalt badhus.",
"##missing_school_or_library##":"Detta hus kan inte utvecklas, eftersom det inte har tillgång till grundläggande utbildningsmöjligheter vare sig från skola eller bibliotek.",
"##missing_barber##":"Detta hus kan inte utvecklas, eftersom det inte har någon lokal tillgång till en barberare.",
"##missing_religion##":"Detta hus kan inte utvecklas, eftersom det inte har tillgång till några lokala möjligheter till religionsutövning.",
"##missing_fountain##":"Detta hus kan inte utvecklas, eftersom det inte har tillgång till ren vattentillförsel från en fontän.",
"##missing_doctor_or_hospital##":"Detta hus kan inte utvecklas, eftersom det i stort sett saknar tillgång till sjukvård. Det saknar tillgång till både klinik och sjukhus.",
"##missing_entertainment_need_more##":"Detta hus kan inte utvecklas, eftersom det visserligen finns god underhållning i området, men inte tillräckligt varierat utbud.",
"##missing_second_wine##":"Detta hus kan inte utvecklas. Det krävs en vinsort till för att tillfredsställa de sysslolösa patriciernas dekadenta livsstil. Öppna en ny handelsväg, eller tillverka ditt eget vin.",
"##missing_wine##":"Detta hus kan inte utvecklas. Det behöver tillgång till vinleveranser från sin lokala marknad innan mer välmående medborgarklasser kommer att flytta in.",
"##missing_oil##":"Detta hus kan inte utvecklas. Det behöver oljeleveranser från sin lokala marknad innan mer välmående medborgarklasser kommer att flytta in.",
"##missing_furniture##":"Detta hus kan inte utvecklas. Det behöver tillgång till möbelleveranser från sin lokala marknad innan mer välmående medborgarklasser kommer att flytta in.",
"##missing_pottery##":"Detta hus kan inte utvecklas. Det behöver leveranser av krukor från sin lokala marknad innan förmögnare medborgarklasser kommer att flytta in.",
"##missing_food_from_market##":"Detta hus kan inte utvecklas. Det har visserligen tillgång till en lokal marknad, men marknaden själv har svårt att få livsmedelsleveranser.",
"##missing_prettyWine_degrade##":"Detta hus kommer snart att förfalla, eftersom staden bara har en enda vinleverantör, och dess krävande invånare klagar över bristande utbud.",
"##missing_furniture_degrade##":"Detta hus kommer snart att förfalla, eftersom det har slut på möbler och dess lokala marknad har ett sporadiskt utbud.",
"##missing_oil_degrade##":"Detta hus kommer snart att förfalla, eftersom det har slut på oljan och dess lokala marknad har ett sporadiskt utbud.",
"##missing_entertainment_degrade##":"Detta hus kommer snart att förfalla, eftersom det knappast finns någon underhållning i området.",
"##missing_entertainment_degrade##":"Detta hus kommer snart att förfalla, eftersom det inte finns tillräckligt med underhållning i området.",
"##missing_doctor_or_hospital_degrade##":"Detta hus kommer snart att förfalla, eftersom det nu har tvivelaktig hälsovård. Det saknas inte bara tillgång till en klinik, utan även tillgången till sjukhus är dålig.",
"##missing_hospital_degrade##":"Detta hus kommer snart att förfalla, eftersom dess tillgång till hälsovård har skurits ned. Tillgången till kliniker är god men det finns inga lokala sjukhus.",
"##missing_wine_degrade##":"Detta hus kommer snart att förfalla, eftersom det har slut på vin och dess lokala marknad har ett sporadiskt utbud.",
"##missing_food_degrade##":"Detta hus kommer snart att förfalla, eftersom det inte har fått några livsmedelsleveranser från en lokal marknad nyligen.",
"##missing_school_or_library_degrade##":"Detta hus kommer snart att förfalla, eftersom det har förlorat alla grundläggande utbildningsmöjligheter från en skola eller ett bibliotek.",
"##missing_religion_degrade##":"Detta hus kommer snart att förfalla, eftersom det har förlorat all tillgång till lokala religiösa byggnader.",
"##missing_bath_degrade##":"Detta hus kommer snart att förfalla, eftersom det har förlorat tillgången till sitt badhus.",
"##missing_barber_degrade##":"Detta hus kommer snart att förfalla, eftersom det har förlorat tillgången till barberare.",
"##missing_third_food_degrade##":"Detta hus kommer snart att förfalla, eftersom det endast har tillgång till 2 typer av livsmedel från sin lokala marknad. Detta avskräcker patricierklasserna.",
"##missing_second_food_degrade##":"Detta hus kommer snart att förfalla, eftersom det endast har tillgång till en enda typ av livsmedel från sin lokala marknad. Detta avskräcker de välbärgade klasserna.",
"##missing_water_degrade##":"Detta hus kommer snart att förfalla, eftersom det saknar tillgång till även den enklaste vattenförsörjning.",
"##missing_fountain_degrade##":"Detta hus kommer snart att förfalla, eftersom det inte har tillgång till rent vatten från en fontän.",
"##missing_pottery_degrade##":"Detta hus kommer snart att förfalla. Det har inte längre tillgång till krukor, och leveranserna till dess lokala marknad är minst sagt opålitliga.",
"##missing_entertainment_amph_degrade##":"Detta hus kommer snart att förfalla. Det finns viss underhållning i området, men inte tillräckligt.",
"##missing_entertainment_also_degrade##":"Detta hus kommer snart att förfalla. Det finns god underhållning i området, men inte tillräckligt varierat utbud.",
"##missing_second_religion_degrade##":"Detta hus kommer snart att förfalla. Dess tillgång till lokala religiösa byggnader har reducerats till endast ett tempel för en enda gud.",
"##missing_library_degrade##":"Detta hus kommer snart att förfalla. Dess tillgång till utbildning har försämrats, eftersom det har förlorat tillgång till sitt bibliotek.",
"##missing_school_degrade##":"Detta hus kommer snart att förfalla. Dess tillgång till utbildning har försämrats, eftersom det har förlorat tillgång till sin skola.",
"##missing_third_religion_degrade##":"Detta hus kommer snart att förfalla. Dess tidigare utmärkta religiösa möjligheter har reducerats, och det har nu endast tillgång till tempel för två gudar.",
"##missing_college_degrade##":"Detta hus kommer snart att förfalla. Dess tidigare utmärkta tillgång till utbildning har försämrats, eftersom det har förlorat tillgången till sin högskola.",
"##low_desirability_degrade##":"Detta hus kommer snart att förfalla. Den sjunkande efterfrågan på boende i detta område drar ner det.",
"##missing_entertainment_colloseum_degrade##":"Detta hus kommer snart att förfalla. Det finns utmärkt underhållning i området, men det är trångt och utbudet är inte tillräckligt varierat för de kräsna patricierna.",
"##missing_food_degrade##":"Detta hus kommer snart att förfalla. Det har visserligen tillgång till en marknad, men marknaden själv har svårt att få livsmedelsleveranser.",
"##missing_market_degrade##":"Detta hus kommer snart att förfalla. Det har förlorat tillgången till en marknad.",
"##missing_doctor__degrade##":"Detta hus kommer snart att förfalla, eftersom dess möjligheter till hälsovård skurits ned. Det finns lokal tillgång till ett sjukhus men det är svårt att hitta en klinik.",
"##hippodrome_no_workers##":"Inget rör sig i hippodromen. Utan arbetare ger den ingen underhållning åt lokalsamhället.",
"##quarry_need_some_workers##":"Detta brott utnyttjar inte maximal kapacitet. Som resultat kommer marmorproduktionen att bli något mindre.",
"##clay_pit_need_some_workers##":"Detta lertag utnyttjar inte full kapacitet. Som resultat kommer lerproduktionen att gå något långsammare.",
"##colloseum_no_workers##":"Detta colosseum är stängt. Utan anställda är det värdelöst som rekreationsanläggning.",
"##trouble_colloseum_have_only_gladiatros##":"Detta colosseum har gladiatorkamp för lokalbefolkningen. Lejon skulle ge mer variation till dödskamperna.",
"##trouble_colloseum_full_work##":"Detta colosseum har både gladiatorkamp och lejonkamper, till lokalsamhällets stora nöje.",
"##trouble_colloseum_have_only_lions##":"Detta colosseum har djurkamp, med lejon från lokala handelsmän. Den skulle också kunna anlita gladiatorer för kamp man mot man.",
"##also_fountain_in_well_area##":"Denna brunn är överflödig för tillfället, eftersom alla hus som den betjänar tar sitt vatten från en fontän.",
"##bridge_extends_city_area##":"Denna bro ger oss mer mark, men ger fri passage både för medborgare och fiender!",
"##oracle_info##":"Orakel ökar efterfrågan på husen i stadsdelen och gör de boende gladare. Denna byggnad tillfredsställer samtliga gudar.",
"##citizen_gods_angry3##":"Den här ståthållaren har ingen respekt för gudarna.",
"##dangerous_crime_risk##":"Detta område är farligt.",
"##extreme_crime_risk##":"Hela detta område är som en jäsande krutdurk! Brottsligheten är epidemisk, och uppror sannolika",
"##reservoir_no_water##":"Denna reservoar fungerar inte eftersom den inte ligger intill vatten eller inte är ansluten till en annan reservoar via akvedukter.",
"##iron_mine_need_some_workers##":"Detta brott utnyttjar inte maximal kapacitet. Malmbrytningen skulle vara mycket effektivare med fler arbetare.",
"##market_no_workers##":"Denna marknad används inte, och levererar inga produkter till lokalsamhället.",
"##market_full_work##":"Denna marknad används",
"##enemies_hard_to_me##":"Denne soldat är för stark för mig!",
"##mopup_formation_text##":"Denna ordning är det effektivaste sättet att hantera resterna av en besegrad armé.",
"##theater_no_have_any_shows##":"Denna teater har sällan några uppsättningar. Den behöver riktiga skådespelare för att kunna erbjuda underhållning.",
"##theater_no_workers##":"Vinden är det enda som rör sig i denna teater. Utan arbetare erbjuder den inga pjäser till lokalbefolkningen.",
"##water_srvc_well##":"Detta område har tillgång till dricksvatten",
"##water_srvc_reservoir##":"Detta område har tillgång till en reservoar via rörledning, vilket gör att fontäner och badhus fungerar",
"##need_reservoir_for_work##":"Denna fontän fungerar inte eftersom den inte ligger i ett område som täcks av rörledningar från en fungerande reservoar.",
"##fountain_not_work##":"Denna fontän fungerar inte eftersom det inte finns tillräckligt med arbetare för att driva den.",
"##fort_has_been_cursed_by_mars##":"Detta fort har förbannats av Mars. Det kommer att dröja innan några soldater vågar sig tillbaka hit.",
"##tarentum_win_text##":"Etruskerna kommer inte att hota Tarentum igen. Bra gjort! Det är sällsynt med en ståthållare som finner rätt balans mellan stadsbyggnation och strid. Låt se om du kan göra om din bravad eller om det bara handlade om tur.",
"##wn_etruscan_soldier##":"En etruskisk soldat",
"##effciency##":"Effektivitet",
"##gmsndwnd_ambient_sound##":"Ljudeffekter",
"##south##":"Syd",
"##southEast##":"Sydost",
"##southWest##":"Sydväst",
"##prefect_gods_angry##":"Jag är rädd för att gudarna kommer att förbanna staden.",
"##legionary_average_life##":"Jag slåss intill döden! Staden är trygg så länge jag lever!",
"##teacher_average_life##":"Jag ger staden åtta av tio poäng.",
"##merchant_notbad_city##":"Jag har kappkört i många värre städer än den här.",
"##cartPusher_cantfind_destination##":"Det skulle gå snabbare att dra varorna till Rom än dit jag ska.",
"##engineer_building_allok##":"Jag behövs knappast. Dessa byggnader är i utmärkt skick.",
"##immigrant_where_my_home##":"Jag är ny i staden. Vet du var man kan få tag i en bostad?",
"##emperor_wrath_by_debt_text##":"Jag är mycket missnöjd. Trots alla pengar jag har investerat i din stad och senatens generösa krediter, har du svikit mig. Din stad har inte betalat tillbaka sina lån. Mitt förtroende för dig var missriktat och jag tvingas nu finna en annan ståthållare i ditt ställe. Du kanske passar bättre i den nya position jag har i åtanke för dig...",
"##landmerchant_good_deals##":"Jag älskar att komma hit. Affärerna går mycket bra.",
"##recruter_low_entertainment##":"Jag arbetar hårt och jag vill roa mig ofta. Men det går inte här. Det finns inget att göra!",
"##cartPusher_gods_angry##":"...religiös, men inte ens jag skulle behandla gudarna på det här sättet.",
"##marketBuyer_need_workers##":"Jag har aldrig sett så många byggnader som behöver fler arbetare.",
"##citizen_high_workless4##":"Jag har aldrig sett så många arbetslösa medborgare förut.",
"##marketBuyer_find_goods##":"Jag ska hämta nya varor.",
"##actor_so_hungry##":"Jag kan inte uppträda utan mer mat.",
"##romeGuard_good_live##":"Jag må vara en simpel soldat, men även jag kan se vilken storslagen stad detta är.",
"##actor_low_entertainment##":"Jag arbetar så hårt jag förmår, men underhållningen i staden räcker inte till på långa vägar.",
"##immigrant_want_to_be_liontamer##":"Jag har hört att det finns arbete här. Jag vill bli lejontämjare.",
"##gladiator_so_hungry##":"Jag är så hungrig att jag kan äta ett lejon!",
"##wt_missioner_normal_life##":"Jag är så glad att vara romare. Du skulle se vad dessa barbarer håller på med i sina hyddor!",
"##teacher_need_workers##":"Otroligt att det finns så många arbetstillfällen här.",
"##scholar_so_hungry##":"Jag svälter ihjäl!",
"##month_1_short##":"Jan",
"##build_senate_for_advisors##":"Bygg senatorbyggnad",
"##click_on_city_for_info_tlp##":"Tryck på stad för information",
}